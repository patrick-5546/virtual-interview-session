module dct_quantization(input logic [7:0][7:0][31:0] mcu, output logic [7:0][7:0][31:0] dct);
	wire[63:0] cos00_term = ((mcu[0][0] * 32'h100) >> 8) + ((mcu[0][1] * 32'h100) >> 8) + ((mcu[0][2] * 32'h100) >> 8) + ((mcu[0][3] * 32'h100) >> 8) + ((mcu[0][4] * 32'h100) >> 8) + ((mcu[0][5] * 32'h100) >> 8) + ((mcu[0][6] * 32'h100) >> 8) + ((mcu[0][7] * 32'h100) >> 8) + ((mcu[1][0] * 32'h100) >> 8) + ((mcu[1][1] * 32'h100) >> 8) + ((mcu[1][2] * 32'h100) >> 8) + ((mcu[1][3] * 32'h100) >> 8) + ((mcu[1][4] * 32'h100) >> 8) + ((mcu[1][5] * 32'h100) >> 8) + ((mcu[1][6] * 32'h100) >> 8) + ((mcu[1][7] * 32'h100) >> 8) + ((mcu[2][0] * 32'h100) >> 8) + ((mcu[2][1] * 32'h100) >> 8) + ((mcu[2][2] * 32'h100) >> 8) + ((mcu[2][3] * 32'h100) >> 8) + ((mcu[2][4] * 32'h100) >> 8) + ((mcu[2][5] * 32'h100) >> 8) + ((mcu[2][6] * 32'h100) >> 8) + ((mcu[2][7] * 32'h100) >> 8) + ((mcu[3][0] * 32'h100) >> 8) + ((mcu[3][1] * 32'h100) >> 8) + ((mcu[3][2] * 32'h100) >> 8) + ((mcu[3][3] * 32'h100) >> 8) + ((mcu[3][4] * 32'h100) >> 8) + ((mcu[3][5] * 32'h100) >> 8) + ((mcu[3][6] * 32'h100) >> 8) + ((mcu[3][7] * 32'h100) >> 8) + ((mcu[4][0] * 32'h100) >> 8) + ((mcu[4][1] * 32'h100) >> 8) + ((mcu[4][2] * 32'h100) >> 8) + ((mcu[4][3] * 32'h100) >> 8) + ((mcu[4][4] * 32'h100) >> 8) + ((mcu[4][5] * 32'h100) >> 8) + ((mcu[4][6] * 32'h100) >> 8) + ((mcu[4][7] * 32'h100) >> 8) + ((mcu[5][0] * 32'h100) >> 8) + ((mcu[5][1] * 32'h100) >> 8) + ((mcu[5][2] * 32'h100) >> 8) + ((mcu[5][3] * 32'h100) >> 8) + ((mcu[5][4] * 32'h100) >> 8) + ((mcu[5][5] * 32'h100) >> 8) + ((mcu[5][6] * 32'h100) >> 8) + ((mcu[5][7] * 32'h100) >> 8) + ((mcu[6][0] * 32'h100) >> 8) + ((mcu[6][1] * 32'h100) >> 8) + ((mcu[6][2] * 32'h100) >> 8) + ((mcu[6][3] * 32'h100) >> 8) + ((mcu[6][4] * 32'h100) >> 8) + ((mcu[6][5] * 32'h100) >> 8) + ((mcu[6][6] * 32'h100) >> 8) + ((mcu[6][7] * 32'h100) >> 8) + ((mcu[7][0] * 32'h100) >> 8) + ((mcu[7][1] * 32'h100) >> 8) + ((mcu[7][2] * 32'h100) >> 8) + ((mcu[7][3] * 32'h100) >> 8) + ((mcu[7][4] * 32'h100) >> 8) + ((mcu[7][5] * 32'h100) >> 8) + ((mcu[7][6] * 32'h100) >> 8) + ((mcu[7][7] * 32'h100) >> 8);
	wire[63:0] cos01_term = ((mcu[0][0] * 32'h0fb) >> 8) + ((mcu[0][1] * 32'h0d4) >> 8) + ((mcu[0][2] * 32'h08e) >> 8) + ((mcu[0][3] * 32'h031) >> 8) + ((mcu[0][4] * -32'h031) >> 8) + ((mcu[0][5] * -32'h08e) >> 8) + ((mcu[0][6] * -32'h0d4) >> 8) + ((mcu[0][7] * -32'h0fb) >> 8) + ((mcu[1][0] * 32'h0fb) >> 8) + ((mcu[1][1] * 32'h0d4) >> 8) + ((mcu[1][2] * 32'h08e) >> 8) + ((mcu[1][3] * 32'h031) >> 8) + ((mcu[1][4] * -32'h031) >> 8) + ((mcu[1][5] * -32'h08e) >> 8) + ((mcu[1][6] * -32'h0d4) >> 8) + ((mcu[1][7] * -32'h0fb) >> 8) + ((mcu[2][0] * 32'h0fb) >> 8) + ((mcu[2][1] * 32'h0d4) >> 8) + ((mcu[2][2] * 32'h08e) >> 8) + ((mcu[2][3] * 32'h031) >> 8) + ((mcu[2][4] * -32'h031) >> 8) + ((mcu[2][5] * -32'h08e) >> 8) + ((mcu[2][6] * -32'h0d4) >> 8) + ((mcu[2][7] * -32'h0fb) >> 8) + ((mcu[3][0] * 32'h0fb) >> 8) + ((mcu[3][1] * 32'h0d4) >> 8) + ((mcu[3][2] * 32'h08e) >> 8) + ((mcu[3][3] * 32'h031) >> 8) + ((mcu[3][4] * -32'h031) >> 8) + ((mcu[3][5] * -32'h08e) >> 8) + ((mcu[3][6] * -32'h0d4) >> 8) + ((mcu[3][7] * -32'h0fb) >> 8) + ((mcu[4][0] * 32'h0fb) >> 8) + ((mcu[4][1] * 32'h0d4) >> 8) + ((mcu[4][2] * 32'h08e) >> 8) + ((mcu[4][3] * 32'h031) >> 8) + ((mcu[4][4] * -32'h031) >> 8) + ((mcu[4][5] * -32'h08e) >> 8) + ((mcu[4][6] * -32'h0d4) >> 8) + ((mcu[4][7] * -32'h0fb) >> 8) + ((mcu[5][0] * 32'h0fb) >> 8) + ((mcu[5][1] * 32'h0d4) >> 8) + ((mcu[5][2] * 32'h08e) >> 8) + ((mcu[5][3] * 32'h031) >> 8) + ((mcu[5][4] * -32'h031) >> 8) + ((mcu[5][5] * -32'h08e) >> 8) + ((mcu[5][6] * -32'h0d4) >> 8) + ((mcu[5][7] * -32'h0fb) >> 8) + ((mcu[6][0] * 32'h0fb) >> 8) + ((mcu[6][1] * 32'h0d4) >> 8) + ((mcu[6][2] * 32'h08e) >> 8) + ((mcu[6][3] * 32'h031) >> 8) + ((mcu[6][4] * -32'h031) >> 8) + ((mcu[6][5] * -32'h08e) >> 8) + ((mcu[6][6] * -32'h0d4) >> 8) + ((mcu[6][7] * -32'h0fb) >> 8) + ((mcu[7][0] * 32'h0fb) >> 8) + ((mcu[7][1] * 32'h0d4) >> 8) + ((mcu[7][2] * 32'h08e) >> 8) + ((mcu[7][3] * 32'h031) >> 8) + ((mcu[7][4] * -32'h031) >> 8) + ((mcu[7][5] * -32'h08e) >> 8) + ((mcu[7][6] * -32'h0d4) >> 8) + ((mcu[7][7] * -32'h0fb) >> 8);
	wire[63:0] cos02_term = ((mcu[0][0] * 32'h0ec) >> 8) + ((mcu[0][1] * 32'h062) >> 8) + ((mcu[0][2] * -32'h062) >> 8) + ((mcu[0][3] * -32'h0ec) >> 8) + ((mcu[0][4] * -32'h0ec) >> 8) + ((mcu[0][5] * -32'h062) >> 8) + ((mcu[0][6] * 32'h062) >> 8) + ((mcu[0][7] * 32'h0ec) >> 8) + ((mcu[1][0] * 32'h0ec) >> 8) + ((mcu[1][1] * 32'h062) >> 8) + ((mcu[1][2] * -32'h062) >> 8) + ((mcu[1][3] * -32'h0ec) >> 8) + ((mcu[1][4] * -32'h0ec) >> 8) + ((mcu[1][5] * -32'h062) >> 8) + ((mcu[1][6] * 32'h062) >> 8) + ((mcu[1][7] * 32'h0ec) >> 8) + ((mcu[2][0] * 32'h0ec) >> 8) + ((mcu[2][1] * 32'h062) >> 8) + ((mcu[2][2] * -32'h062) >> 8) + ((mcu[2][3] * -32'h0ec) >> 8) + ((mcu[2][4] * -32'h0ec) >> 8) + ((mcu[2][5] * -32'h062) >> 8) + ((mcu[2][6] * 32'h062) >> 8) + ((mcu[2][7] * 32'h0ec) >> 8) + ((mcu[3][0] * 32'h0ec) >> 8) + ((mcu[3][1] * 32'h062) >> 8) + ((mcu[3][2] * -32'h062) >> 8) + ((mcu[3][3] * -32'h0ec) >> 8) + ((mcu[3][4] * -32'h0ec) >> 8) + ((mcu[3][5] * -32'h062) >> 8) + ((mcu[3][6] * 32'h062) >> 8) + ((mcu[3][7] * 32'h0ec) >> 8) + ((mcu[4][0] * 32'h0ec) >> 8) + ((mcu[4][1] * 32'h062) >> 8) + ((mcu[4][2] * -32'h062) >> 8) + ((mcu[4][3] * -32'h0ec) >> 8) + ((mcu[4][4] * -32'h0ec) >> 8) + ((mcu[4][5] * -32'h062) >> 8) + ((mcu[4][6] * 32'h062) >> 8) + ((mcu[4][7] * 32'h0ec) >> 8) + ((mcu[5][0] * 32'h0ec) >> 8) + ((mcu[5][1] * 32'h062) >> 8) + ((mcu[5][2] * -32'h062) >> 8) + ((mcu[5][3] * -32'h0ec) >> 8) + ((mcu[5][4] * -32'h0ec) >> 8) + ((mcu[5][5] * -32'h062) >> 8) + ((mcu[5][6] * 32'h062) >> 8) + ((mcu[5][7] * 32'h0ec) >> 8) + ((mcu[6][0] * 32'h0ec) >> 8) + ((mcu[6][1] * 32'h062) >> 8) + ((mcu[6][2] * -32'h062) >> 8) + ((mcu[6][3] * -32'h0ec) >> 8) + ((mcu[6][4] * -32'h0ec) >> 8) + ((mcu[6][5] * -32'h062) >> 8) + ((mcu[6][6] * 32'h062) >> 8) + ((mcu[6][7] * 32'h0ec) >> 8) + ((mcu[7][0] * 32'h0ec) >> 8) + ((mcu[7][1] * 32'h062) >> 8) + ((mcu[7][2] * -32'h062) >> 8) + ((mcu[7][3] * -32'h0ec) >> 8) + ((mcu[7][4] * -32'h0ec) >> 8) + ((mcu[7][5] * -32'h062) >> 8) + ((mcu[7][6] * 32'h062) >> 8) + ((mcu[7][7] * 32'h0ec) >> 8);
	wire[63:0] cos03_term = ((mcu[0][0] * 32'h0d4) >> 8) + ((mcu[0][1] * -32'h031) >> 8) + ((mcu[0][2] * -32'h0fb) >> 8) + ((mcu[0][3] * -32'h08e) >> 8) + ((mcu[0][4] * 32'h08e) >> 8) + ((mcu[0][5] * 32'h0fb) >> 8) + ((mcu[0][6] * 32'h031) >> 8) + ((mcu[0][7] * -32'h0d4) >> 8) + ((mcu[1][0] * 32'h0d4) >> 8) + ((mcu[1][1] * -32'h031) >> 8) + ((mcu[1][2] * -32'h0fb) >> 8) + ((mcu[1][3] * -32'h08e) >> 8) + ((mcu[1][4] * 32'h08e) >> 8) + ((mcu[1][5] * 32'h0fb) >> 8) + ((mcu[1][6] * 32'h031) >> 8) + ((mcu[1][7] * -32'h0d4) >> 8) + ((mcu[2][0] * 32'h0d4) >> 8) + ((mcu[2][1] * -32'h031) >> 8) + ((mcu[2][2] * -32'h0fb) >> 8) + ((mcu[2][3] * -32'h08e) >> 8) + ((mcu[2][4] * 32'h08e) >> 8) + ((mcu[2][5] * 32'h0fb) >> 8) + ((mcu[2][6] * 32'h031) >> 8) + ((mcu[2][7] * -32'h0d4) >> 8) + ((mcu[3][0] * 32'h0d4) >> 8) + ((mcu[3][1] * -32'h031) >> 8) + ((mcu[3][2] * -32'h0fb) >> 8) + ((mcu[3][3] * -32'h08e) >> 8) + ((mcu[3][4] * 32'h08e) >> 8) + ((mcu[3][5] * 32'h0fb) >> 8) + ((mcu[3][6] * 32'h031) >> 8) + ((mcu[3][7] * -32'h0d4) >> 8) + ((mcu[4][0] * 32'h0d4) >> 8) + ((mcu[4][1] * -32'h031) >> 8) + ((mcu[4][2] * -32'h0fb) >> 8) + ((mcu[4][3] * -32'h08e) >> 8) + ((mcu[4][4] * 32'h08e) >> 8) + ((mcu[4][5] * 32'h0fb) >> 8) + ((mcu[4][6] * 32'h031) >> 8) + ((mcu[4][7] * -32'h0d4) >> 8) + ((mcu[5][0] * 32'h0d4) >> 8) + ((mcu[5][1] * -32'h031) >> 8) + ((mcu[5][2] * -32'h0fb) >> 8) + ((mcu[5][3] * -32'h08e) >> 8) + ((mcu[5][4] * 32'h08e) >> 8) + ((mcu[5][5] * 32'h0fb) >> 8) + ((mcu[5][6] * 32'h031) >> 8) + ((mcu[5][7] * -32'h0d4) >> 8) + ((mcu[6][0] * 32'h0d4) >> 8) + ((mcu[6][1] * -32'h031) >> 8) + ((mcu[6][2] * -32'h0fb) >> 8) + ((mcu[6][3] * -32'h08e) >> 8) + ((mcu[6][4] * 32'h08e) >> 8) + ((mcu[6][5] * 32'h0fb) >> 8) + ((mcu[6][6] * 32'h031) >> 8) + ((mcu[6][7] * -32'h0d4) >> 8) + ((mcu[7][0] * 32'h0d4) >> 8) + ((mcu[7][1] * -32'h031) >> 8) + ((mcu[7][2] * -32'h0fb) >> 8) + ((mcu[7][3] * -32'h08e) >> 8) + ((mcu[7][4] * 32'h08e) >> 8) + ((mcu[7][5] * 32'h0fb) >> 8) + ((mcu[7][6] * 32'h031) >> 8) + ((mcu[7][7] * -32'h0d4) >> 8);
	wire[63:0] cos04_term = ((mcu[0][0] * 32'h0b4) >> 8) + ((mcu[0][1] * -32'h0b4) >> 8) + ((mcu[0][2] * -32'h0b4) >> 8) + ((mcu[0][3] * 32'h0b4) >> 8) + ((mcu[0][4] * 32'h0b4) >> 8) + ((mcu[0][5] * -32'h0b4) >> 8) + ((mcu[0][6] * -32'h0b4) >> 8) + ((mcu[0][7] * 32'h0b4) >> 8) + ((mcu[1][0] * 32'h0b4) >> 8) + ((mcu[1][1] * -32'h0b4) >> 8) + ((mcu[1][2] * -32'h0b4) >> 8) + ((mcu[1][3] * 32'h0b4) >> 8) + ((mcu[1][4] * 32'h0b4) >> 8) + ((mcu[1][5] * -32'h0b4) >> 8) + ((mcu[1][6] * -32'h0b4) >> 8) + ((mcu[1][7] * 32'h0b4) >> 8) + ((mcu[2][0] * 32'h0b4) >> 8) + ((mcu[2][1] * -32'h0b4) >> 8) + ((mcu[2][2] * -32'h0b4) >> 8) + ((mcu[2][3] * 32'h0b4) >> 8) + ((mcu[2][4] * 32'h0b4) >> 8) + ((mcu[2][5] * -32'h0b4) >> 8) + ((mcu[2][6] * -32'h0b4) >> 8) + ((mcu[2][7] * 32'h0b4) >> 8) + ((mcu[3][0] * 32'h0b4) >> 8) + ((mcu[3][1] * -32'h0b4) >> 8) + ((mcu[3][2] * -32'h0b4) >> 8) + ((mcu[3][3] * 32'h0b4) >> 8) + ((mcu[3][4] * 32'h0b4) >> 8) + ((mcu[3][5] * -32'h0b4) >> 8) + ((mcu[3][6] * -32'h0b4) >> 8) + ((mcu[3][7] * 32'h0b4) >> 8) + ((mcu[4][0] * 32'h0b4) >> 8) + ((mcu[4][1] * -32'h0b4) >> 8) + ((mcu[4][2] * -32'h0b4) >> 8) + ((mcu[4][3] * 32'h0b4) >> 8) + ((mcu[4][4] * 32'h0b4) >> 8) + ((mcu[4][5] * -32'h0b4) >> 8) + ((mcu[4][6] * -32'h0b4) >> 8) + ((mcu[4][7] * 32'h0b4) >> 8) + ((mcu[5][0] * 32'h0b4) >> 8) + ((mcu[5][1] * -32'h0b4) >> 8) + ((mcu[5][2] * -32'h0b4) >> 8) + ((mcu[5][3] * 32'h0b4) >> 8) + ((mcu[5][4] * 32'h0b4) >> 8) + ((mcu[5][5] * -32'h0b4) >> 8) + ((mcu[5][6] * -32'h0b4) >> 8) + ((mcu[5][7] * 32'h0b4) >> 8) + ((mcu[6][0] * 32'h0b4) >> 8) + ((mcu[6][1] * -32'h0b4) >> 8) + ((mcu[6][2] * -32'h0b4) >> 8) + ((mcu[6][3] * 32'h0b4) >> 8) + ((mcu[6][4] * 32'h0b4) >> 8) + ((mcu[6][5] * -32'h0b4) >> 8) + ((mcu[6][6] * -32'h0b4) >> 8) + ((mcu[6][7] * 32'h0b4) >> 8) + ((mcu[7][0] * 32'h0b4) >> 8) + ((mcu[7][1] * -32'h0b4) >> 8) + ((mcu[7][2] * -32'h0b4) >> 8) + ((mcu[7][3] * 32'h0b4) >> 8) + ((mcu[7][4] * 32'h0b4) >> 8) + ((mcu[7][5] * -32'h0b4) >> 8) + ((mcu[7][6] * -32'h0b4) >> 8) + ((mcu[7][7] * 32'h0b4) >> 8);
	wire[63:0] cos05_term = ((mcu[0][0] * 32'h08e) >> 8) + ((mcu[0][1] * -32'h0fb) >> 8) + ((mcu[0][2] * 32'h031) >> 8) + ((mcu[0][3] * 32'h0d4) >> 8) + ((mcu[0][4] * -32'h0d4) >> 8) + ((mcu[0][5] * -32'h031) >> 8) + ((mcu[0][6] * 32'h0fb) >> 8) + ((mcu[0][7] * -32'h08e) >> 8) + ((mcu[1][0] * 32'h08e) >> 8) + ((mcu[1][1] * -32'h0fb) >> 8) + ((mcu[1][2] * 32'h031) >> 8) + ((mcu[1][3] * 32'h0d4) >> 8) + ((mcu[1][4] * -32'h0d4) >> 8) + ((mcu[1][5] * -32'h031) >> 8) + ((mcu[1][6] * 32'h0fb) >> 8) + ((mcu[1][7] * -32'h08e) >> 8) + ((mcu[2][0] * 32'h08e) >> 8) + ((mcu[2][1] * -32'h0fb) >> 8) + ((mcu[2][2] * 32'h031) >> 8) + ((mcu[2][3] * 32'h0d4) >> 8) + ((mcu[2][4] * -32'h0d4) >> 8) + ((mcu[2][5] * -32'h031) >> 8) + ((mcu[2][6] * 32'h0fb) >> 8) + ((mcu[2][7] * -32'h08e) >> 8) + ((mcu[3][0] * 32'h08e) >> 8) + ((mcu[3][1] * -32'h0fb) >> 8) + ((mcu[3][2] * 32'h031) >> 8) + ((mcu[3][3] * 32'h0d4) >> 8) + ((mcu[3][4] * -32'h0d4) >> 8) + ((mcu[3][5] * -32'h031) >> 8) + ((mcu[3][6] * 32'h0fb) >> 8) + ((mcu[3][7] * -32'h08e) >> 8) + ((mcu[4][0] * 32'h08e) >> 8) + ((mcu[4][1] * -32'h0fb) >> 8) + ((mcu[4][2] * 32'h031) >> 8) + ((mcu[4][3] * 32'h0d4) >> 8) + ((mcu[4][4] * -32'h0d4) >> 8) + ((mcu[4][5] * -32'h031) >> 8) + ((mcu[4][6] * 32'h0fb) >> 8) + ((mcu[4][7] * -32'h08e) >> 8) + ((mcu[5][0] * 32'h08e) >> 8) + ((mcu[5][1] * -32'h0fb) >> 8) + ((mcu[5][2] * 32'h031) >> 8) + ((mcu[5][3] * 32'h0d4) >> 8) + ((mcu[5][4] * -32'h0d4) >> 8) + ((mcu[5][5] * -32'h031) >> 8) + ((mcu[5][6] * 32'h0fb) >> 8) + ((mcu[5][7] * -32'h08e) >> 8) + ((mcu[6][0] * 32'h08e) >> 8) + ((mcu[6][1] * -32'h0fb) >> 8) + ((mcu[6][2] * 32'h031) >> 8) + ((mcu[6][3] * 32'h0d4) >> 8) + ((mcu[6][4] * -32'h0d4) >> 8) + ((mcu[6][5] * -32'h031) >> 8) + ((mcu[6][6] * 32'h0fb) >> 8) + ((mcu[6][7] * -32'h08e) >> 8) + ((mcu[7][0] * 32'h08e) >> 8) + ((mcu[7][1] * -32'h0fb) >> 8) + ((mcu[7][2] * 32'h031) >> 8) + ((mcu[7][3] * 32'h0d4) >> 8) + ((mcu[7][4] * -32'h0d4) >> 8) + ((mcu[7][5] * -32'h031) >> 8) + ((mcu[7][6] * 32'h0fb) >> 8) + ((mcu[7][7] * -32'h08e) >> 8);
	wire[63:0] cos06_term = ((mcu[0][0] * 32'h062) >> 8) + ((mcu[0][1] * -32'h0ec) >> 8) + ((mcu[0][2] * 32'h0ec) >> 8) + ((mcu[0][3] * -32'h062) >> 8) + ((mcu[0][4] * -32'h062) >> 8) + ((mcu[0][5] * 32'h0ec) >> 8) + ((mcu[0][6] * -32'h0ec) >> 8) + ((mcu[0][7] * 32'h062) >> 8) + ((mcu[1][0] * 32'h062) >> 8) + ((mcu[1][1] * -32'h0ec) >> 8) + ((mcu[1][2] * 32'h0ec) >> 8) + ((mcu[1][3] * -32'h062) >> 8) + ((mcu[1][4] * -32'h062) >> 8) + ((mcu[1][5] * 32'h0ec) >> 8) + ((mcu[1][6] * -32'h0ec) >> 8) + ((mcu[1][7] * 32'h062) >> 8) + ((mcu[2][0] * 32'h062) >> 8) + ((mcu[2][1] * -32'h0ec) >> 8) + ((mcu[2][2] * 32'h0ec) >> 8) + ((mcu[2][3] * -32'h062) >> 8) + ((mcu[2][4] * -32'h062) >> 8) + ((mcu[2][5] * 32'h0ec) >> 8) + ((mcu[2][6] * -32'h0ec) >> 8) + ((mcu[2][7] * 32'h062) >> 8) + ((mcu[3][0] * 32'h062) >> 8) + ((mcu[3][1] * -32'h0ec) >> 8) + ((mcu[3][2] * 32'h0ec) >> 8) + ((mcu[3][3] * -32'h062) >> 8) + ((mcu[3][4] * -32'h062) >> 8) + ((mcu[3][5] * 32'h0ec) >> 8) + ((mcu[3][6] * -32'h0ec) >> 8) + ((mcu[3][7] * 32'h062) >> 8) + ((mcu[4][0] * 32'h062) >> 8) + ((mcu[4][1] * -32'h0ec) >> 8) + ((mcu[4][2] * 32'h0ec) >> 8) + ((mcu[4][3] * -32'h062) >> 8) + ((mcu[4][4] * -32'h062) >> 8) + ((mcu[4][5] * 32'h0ec) >> 8) + ((mcu[4][6] * -32'h0ec) >> 8) + ((mcu[4][7] * 32'h062) >> 8) + ((mcu[5][0] * 32'h062) >> 8) + ((mcu[5][1] * -32'h0ec) >> 8) + ((mcu[5][2] * 32'h0ec) >> 8) + ((mcu[5][3] * -32'h062) >> 8) + ((mcu[5][4] * -32'h062) >> 8) + ((mcu[5][5] * 32'h0ec) >> 8) + ((mcu[5][6] * -32'h0ec) >> 8) + ((mcu[5][7] * 32'h062) >> 8) + ((mcu[6][0] * 32'h062) >> 8) + ((mcu[6][1] * -32'h0ec) >> 8) + ((mcu[6][2] * 32'h0ec) >> 8) + ((mcu[6][3] * -32'h062) >> 8) + ((mcu[6][4] * -32'h062) >> 8) + ((mcu[6][5] * 32'h0ec) >> 8) + ((mcu[6][6] * -32'h0ec) >> 8) + ((mcu[6][7] * 32'h062) >> 8) + ((mcu[7][0] * 32'h062) >> 8) + ((mcu[7][1] * -32'h0ec) >> 8) + ((mcu[7][2] * 32'h0ec) >> 8) + ((mcu[7][3] * -32'h062) >> 8) + ((mcu[7][4] * -32'h062) >> 8) + ((mcu[7][5] * 32'h0ec) >> 8) + ((mcu[7][6] * -32'h0ec) >> 8) + ((mcu[7][7] * 32'h062) >> 8);
	wire[63:0] cos07_term = ((mcu[0][0] * 32'h031) >> 8) + ((mcu[0][1] * -32'h08e) >> 8) + ((mcu[0][2] * 32'h0d4) >> 8) + ((mcu[0][3] * -32'h0fb) >> 8) + ((mcu[0][4] * 32'h0fb) >> 8) + ((mcu[0][5] * -32'h0d4) >> 8) + ((mcu[0][6] * 32'h08e) >> 8) + ((mcu[0][7] * -32'h031) >> 8) + ((mcu[1][0] * 32'h031) >> 8) + ((mcu[1][1] * -32'h08e) >> 8) + ((mcu[1][2] * 32'h0d4) >> 8) + ((mcu[1][3] * -32'h0fb) >> 8) + ((mcu[1][4] * 32'h0fb) >> 8) + ((mcu[1][5] * -32'h0d4) >> 8) + ((mcu[1][6] * 32'h08e) >> 8) + ((mcu[1][7] * -32'h031) >> 8) + ((mcu[2][0] * 32'h031) >> 8) + ((mcu[2][1] * -32'h08e) >> 8) + ((mcu[2][2] * 32'h0d4) >> 8) + ((mcu[2][3] * -32'h0fb) >> 8) + ((mcu[2][4] * 32'h0fb) >> 8) + ((mcu[2][5] * -32'h0d4) >> 8) + ((mcu[2][6] * 32'h08e) >> 8) + ((mcu[2][7] * -32'h031) >> 8) + ((mcu[3][0] * 32'h031) >> 8) + ((mcu[3][1] * -32'h08e) >> 8) + ((mcu[3][2] * 32'h0d4) >> 8) + ((mcu[3][3] * -32'h0fb) >> 8) + ((mcu[3][4] * 32'h0fb) >> 8) + ((mcu[3][5] * -32'h0d4) >> 8) + ((mcu[3][6] * 32'h08e) >> 8) + ((mcu[3][7] * -32'h031) >> 8) + ((mcu[4][0] * 32'h031) >> 8) + ((mcu[4][1] * -32'h08e) >> 8) + ((mcu[4][2] * 32'h0d4) >> 8) + ((mcu[4][3] * -32'h0fb) >> 8) + ((mcu[4][4] * 32'h0fb) >> 8) + ((mcu[4][5] * -32'h0d4) >> 8) + ((mcu[4][6] * 32'h08e) >> 8) + ((mcu[4][7] * -32'h031) >> 8) + ((mcu[5][0] * 32'h031) >> 8) + ((mcu[5][1] * -32'h08e) >> 8) + ((mcu[5][2] * 32'h0d4) >> 8) + ((mcu[5][3] * -32'h0fb) >> 8) + ((mcu[5][4] * 32'h0fb) >> 8) + ((mcu[5][5] * -32'h0d4) >> 8) + ((mcu[5][6] * 32'h08e) >> 8) + ((mcu[5][7] * -32'h031) >> 8) + ((mcu[6][0] * 32'h031) >> 8) + ((mcu[6][1] * -32'h08e) >> 8) + ((mcu[6][2] * 32'h0d4) >> 8) + ((mcu[6][3] * -32'h0fb) >> 8) + ((mcu[6][4] * 32'h0fb) >> 8) + ((mcu[6][5] * -32'h0d4) >> 8) + ((mcu[6][6] * 32'h08e) >> 8) + ((mcu[6][7] * -32'h031) >> 8) + ((mcu[7][0] * 32'h031) >> 8) + ((mcu[7][1] * -32'h08e) >> 8) + ((mcu[7][2] * 32'h0d4) >> 8) + ((mcu[7][3] * -32'h0fb) >> 8) + ((mcu[7][4] * 32'h0fb) >> 8) + ((mcu[7][5] * -32'h0d4) >> 8) + ((mcu[7][6] * 32'h08e) >> 8) + ((mcu[7][7] * -32'h031) >> 8);
	wire[63:0] cos10_term = ((mcu[0][0] * 32'h0fb) >> 8) + ((mcu[0][1] * 32'h0fb) >> 8) + ((mcu[0][2] * 32'h0fb) >> 8) + ((mcu[0][3] * 32'h0fb) >> 8) + ((mcu[0][4] * 32'h0fb) >> 8) + ((mcu[0][5] * 32'h0fb) >> 8) + ((mcu[0][6] * 32'h0fb) >> 8) + ((mcu[0][7] * 32'h0fb) >> 8) + ((mcu[1][0] * 32'h0d4) >> 8) + ((mcu[1][1] * 32'h0d4) >> 8) + ((mcu[1][2] * 32'h0d4) >> 8) + ((mcu[1][3] * 32'h0d4) >> 8) + ((mcu[1][4] * 32'h0d4) >> 8) + ((mcu[1][5] * 32'h0d4) >> 8) + ((mcu[1][6] * 32'h0d4) >> 8) + ((mcu[1][7] * 32'h0d4) >> 8) + ((mcu[2][0] * 32'h08e) >> 8) + ((mcu[2][1] * 32'h08e) >> 8) + ((mcu[2][2] * 32'h08e) >> 8) + ((mcu[2][3] * 32'h08e) >> 8) + ((mcu[2][4] * 32'h08e) >> 8) + ((mcu[2][5] * 32'h08e) >> 8) + ((mcu[2][6] * 32'h08e) >> 8) + ((mcu[2][7] * 32'h08e) >> 8) + ((mcu[3][0] * 32'h031) >> 8) + ((mcu[3][1] * 32'h031) >> 8) + ((mcu[3][2] * 32'h031) >> 8) + ((mcu[3][3] * 32'h031) >> 8) + ((mcu[3][4] * 32'h031) >> 8) + ((mcu[3][5] * 32'h031) >> 8) + ((mcu[3][6] * 32'h031) >> 8) + ((mcu[3][7] * 32'h031) >> 8) + ((mcu[4][0] * -32'h031) >> 8) + ((mcu[4][1] * -32'h031) >> 8) + ((mcu[4][2] * -32'h031) >> 8) + ((mcu[4][3] * -32'h031) >> 8) + ((mcu[4][4] * -32'h031) >> 8) + ((mcu[4][5] * -32'h031) >> 8) + ((mcu[4][6] * -32'h031) >> 8) + ((mcu[4][7] * -32'h031) >> 8) + ((mcu[5][0] * -32'h08e) >> 8) + ((mcu[5][1] * -32'h08e) >> 8) + ((mcu[5][2] * -32'h08e) >> 8) + ((mcu[5][3] * -32'h08e) >> 8) + ((mcu[5][4] * -32'h08e) >> 8) + ((mcu[5][5] * -32'h08e) >> 8) + ((mcu[5][6] * -32'h08e) >> 8) + ((mcu[5][7] * -32'h08e) >> 8) + ((mcu[6][0] * -32'h0d4) >> 8) + ((mcu[6][1] * -32'h0d4) >> 8) + ((mcu[6][2] * -32'h0d4) >> 8) + ((mcu[6][3] * -32'h0d4) >> 8) + ((mcu[6][4] * -32'h0d4) >> 8) + ((mcu[6][5] * -32'h0d4) >> 8) + ((mcu[6][6] * -32'h0d4) >> 8) + ((mcu[6][7] * -32'h0d4) >> 8) + ((mcu[7][0] * -32'h0fb) >> 8) + ((mcu[7][1] * -32'h0fb) >> 8) + ((mcu[7][2] * -32'h0fb) >> 8) + ((mcu[7][3] * -32'h0fb) >> 8) + ((mcu[7][4] * -32'h0fb) >> 8) + ((mcu[7][5] * -32'h0fb) >> 8) + ((mcu[7][6] * -32'h0fb) >> 8) + ((mcu[7][7] * -32'h0fb) >> 8);
	wire[63:0] cos11_term = ((mcu[0][0] * 32'h0f6) >> 8) + ((mcu[0][1] * 32'h0d0) >> 8) + ((mcu[0][2] * 32'h08b) >> 8) + ((mcu[0][3] * 32'h030) >> 8) + ((mcu[0][4] * -32'h030) >> 8) + ((mcu[0][5] * -32'h08b) >> 8) + ((mcu[0][6] * -32'h0d0) >> 8) + ((mcu[0][7] * -32'h0f6) >> 8) + ((mcu[1][0] * 32'h0d0) >> 8) + ((mcu[1][1] * 32'h0b0) >> 8) + ((mcu[1][2] * 32'h076) >> 8) + ((mcu[1][3] * 32'h029) >> 8) + ((mcu[1][4] * -32'h029) >> 8) + ((mcu[1][5] * -32'h076) >> 8) + ((mcu[1][6] * -32'h0b0) >> 8) + ((mcu[1][7] * -32'h0d0) >> 8) + ((mcu[2][0] * 32'h08b) >> 8) + ((mcu[2][1] * 32'h076) >> 8) + ((mcu[2][2] * 32'h04f) >> 8) + ((mcu[2][3] * 32'h01b) >> 8) + ((mcu[2][4] * -32'h01b) >> 8) + ((mcu[2][5] * -32'h04f) >> 8) + ((mcu[2][6] * -32'h076) >> 8) + ((mcu[2][7] * -32'h08b) >> 8) + ((mcu[3][0] * 32'h030) >> 8) + ((mcu[3][1] * 32'h029) >> 8) + ((mcu[3][2] * 32'h01b) >> 8) + ((mcu[3][3] * 32'h009) >> 8) + ((mcu[3][4] * -32'h009) >> 8) + ((mcu[3][5] * -32'h01b) >> 8) + ((mcu[3][6] * -32'h029) >> 8) + ((mcu[3][7] * -32'h030) >> 8) + ((mcu[4][0] * -32'h030) >> 8) + ((mcu[4][1] * -32'h029) >> 8) + ((mcu[4][2] * -32'h01b) >> 8) + ((mcu[4][3] * -32'h009) >> 8) + ((mcu[4][4] * 32'h009) >> 8) + ((mcu[4][5] * 32'h01b) >> 8) + ((mcu[4][6] * 32'h029) >> 8) + ((mcu[4][7] * 32'h030) >> 8) + ((mcu[5][0] * -32'h08b) >> 8) + ((mcu[5][1] * -32'h076) >> 8) + ((mcu[5][2] * -32'h04f) >> 8) + ((mcu[5][3] * -32'h01b) >> 8) + ((mcu[5][4] * 32'h01b) >> 8) + ((mcu[5][5] * 32'h04f) >> 8) + ((mcu[5][6] * 32'h076) >> 8) + ((mcu[5][7] * 32'h08b) >> 8) + ((mcu[6][0] * -32'h0d0) >> 8) + ((mcu[6][1] * -32'h0b0) >> 8) + ((mcu[6][2] * -32'h076) >> 8) + ((mcu[6][3] * -32'h029) >> 8) + ((mcu[6][4] * 32'h029) >> 8) + ((mcu[6][5] * 32'h076) >> 8) + ((mcu[6][6] * 32'h0b0) >> 8) + ((mcu[6][7] * 32'h0d0) >> 8) + ((mcu[7][0] * -32'h0f6) >> 8) + ((mcu[7][1] * -32'h0d0) >> 8) + ((mcu[7][2] * -32'h08b) >> 8) + ((mcu[7][3] * -32'h030) >> 8) + ((mcu[7][4] * 32'h030) >> 8) + ((mcu[7][5] * 32'h08b) >> 8) + ((mcu[7][6] * 32'h0d0) >> 8) + ((mcu[7][7] * 32'h0f6) >> 8);
	wire[63:0] cos12_term = ((mcu[0][0] * 32'h0e7) >> 8) + ((mcu[0][1] * 32'h060) >> 8) + ((mcu[0][2] * -32'h060) >> 8) + ((mcu[0][3] * -32'h0e7) >> 8) + ((mcu[0][4] * -32'h0e7) >> 8) + ((mcu[0][5] * -32'h060) >> 8) + ((mcu[0][6] * 32'h060) >> 8) + ((mcu[0][7] * 32'h0e7) >> 8) + ((mcu[1][0] * 32'h0c4) >> 8) + ((mcu[1][1] * 32'h051) >> 8) + ((mcu[1][2] * -32'h051) >> 8) + ((mcu[1][3] * -32'h0c4) >> 8) + ((mcu[1][4] * -32'h0c4) >> 8) + ((mcu[1][5] * -32'h051) >> 8) + ((mcu[1][6] * 32'h051) >> 8) + ((mcu[1][7] * 32'h0c4) >> 8) + ((mcu[2][0] * 32'h083) >> 8) + ((mcu[2][1] * 32'h036) >> 8) + ((mcu[2][2] * -32'h036) >> 8) + ((mcu[2][3] * -32'h083) >> 8) + ((mcu[2][4] * -32'h083) >> 8) + ((mcu[2][5] * -32'h036) >> 8) + ((mcu[2][6] * 32'h036) >> 8) + ((mcu[2][7] * 32'h083) >> 8) + ((mcu[3][0] * 32'h02e) >> 8) + ((mcu[3][1] * 32'h013) >> 8) + ((mcu[3][2] * -32'h013) >> 8) + ((mcu[3][3] * -32'h02e) >> 8) + ((mcu[3][4] * -32'h02e) >> 8) + ((mcu[3][5] * -32'h013) >> 8) + ((mcu[3][6] * 32'h013) >> 8) + ((mcu[3][7] * 32'h02e) >> 8) + ((mcu[4][0] * -32'h02e) >> 8) + ((mcu[4][1] * -32'h013) >> 8) + ((mcu[4][2] * 32'h013) >> 8) + ((mcu[4][3] * 32'h02e) >> 8) + ((mcu[4][4] * 32'h02e) >> 8) + ((mcu[4][5] * 32'h013) >> 8) + ((mcu[4][6] * -32'h013) >> 8) + ((mcu[4][7] * -32'h02e) >> 8) + ((mcu[5][0] * -32'h083) >> 8) + ((mcu[5][1] * -32'h036) >> 8) + ((mcu[5][2] * 32'h036) >> 8) + ((mcu[5][3] * 32'h083) >> 8) + ((mcu[5][4] * 32'h083) >> 8) + ((mcu[5][5] * 32'h036) >> 8) + ((mcu[5][6] * -32'h036) >> 8) + ((mcu[5][7] * -32'h083) >> 8) + ((mcu[6][0] * -32'h0c4) >> 8) + ((mcu[6][1] * -32'h051) >> 8) + ((mcu[6][2] * 32'h051) >> 8) + ((mcu[6][3] * 32'h0c4) >> 8) + ((mcu[6][4] * 32'h0c4) >> 8) + ((mcu[6][5] * 32'h051) >> 8) + ((mcu[6][6] * -32'h051) >> 8) + ((mcu[6][7] * -32'h0c4) >> 8) + ((mcu[7][0] * -32'h0e7) >> 8) + ((mcu[7][1] * -32'h060) >> 8) + ((mcu[7][2] * 32'h060) >> 8) + ((mcu[7][3] * 32'h0e7) >> 8) + ((mcu[7][4] * 32'h0e7) >> 8) + ((mcu[7][5] * 32'h060) >> 8) + ((mcu[7][6] * -32'h060) >> 8) + ((mcu[7][7] * -32'h0e7) >> 8);
	wire[63:0] cos13_term = ((mcu[0][0] * 32'h0d0) >> 8) + ((mcu[0][1] * -32'h030) >> 8) + ((mcu[0][2] * -32'h0f6) >> 8) + ((mcu[0][3] * -32'h08b) >> 8) + ((mcu[0][4] * 32'h08b) >> 8) + ((mcu[0][5] * 32'h0f6) >> 8) + ((mcu[0][6] * 32'h030) >> 8) + ((mcu[0][7] * -32'h0d0) >> 8) + ((mcu[1][0] * 32'h0b0) >> 8) + ((mcu[1][1] * -32'h029) >> 8) + ((mcu[1][2] * -32'h0d0) >> 8) + ((mcu[1][3] * -32'h076) >> 8) + ((mcu[1][4] * 32'h076) >> 8) + ((mcu[1][5] * 32'h0d0) >> 8) + ((mcu[1][6] * 32'h029) >> 8) + ((mcu[1][7] * -32'h0b0) >> 8) + ((mcu[2][0] * 32'h076) >> 8) + ((mcu[2][1] * -32'h01b) >> 8) + ((mcu[2][2] * -32'h08b) >> 8) + ((mcu[2][3] * -32'h04f) >> 8) + ((mcu[2][4] * 32'h04f) >> 8) + ((mcu[2][5] * 32'h08b) >> 8) + ((mcu[2][6] * 32'h01b) >> 8) + ((mcu[2][7] * -32'h076) >> 8) + ((mcu[3][0] * 32'h029) >> 8) + ((mcu[3][1] * -32'h009) >> 8) + ((mcu[3][2] * -32'h030) >> 8) + ((mcu[3][3] * -32'h01b) >> 8) + ((mcu[3][4] * 32'h01b) >> 8) + ((mcu[3][5] * 32'h030) >> 8) + ((mcu[3][6] * 32'h009) >> 8) + ((mcu[3][7] * -32'h029) >> 8) + ((mcu[4][0] * -32'h029) >> 8) + ((mcu[4][1] * 32'h009) >> 8) + ((mcu[4][2] * 32'h030) >> 8) + ((mcu[4][3] * 32'h01b) >> 8) + ((mcu[4][4] * -32'h01b) >> 8) + ((mcu[4][5] * -32'h030) >> 8) + ((mcu[4][6] * -32'h009) >> 8) + ((mcu[4][7] * 32'h029) >> 8) + ((mcu[5][0] * -32'h076) >> 8) + ((mcu[5][1] * 32'h01b) >> 8) + ((mcu[5][2] * 32'h08b) >> 8) + ((mcu[5][3] * 32'h04f) >> 8) + ((mcu[5][4] * -32'h04f) >> 8) + ((mcu[5][5] * -32'h08b) >> 8) + ((mcu[5][6] * -32'h01b) >> 8) + ((mcu[5][7] * 32'h076) >> 8) + ((mcu[6][0] * -32'h0b0) >> 8) + ((mcu[6][1] * 32'h029) >> 8) + ((mcu[6][2] * 32'h0d0) >> 8) + ((mcu[6][3] * 32'h076) >> 8) + ((mcu[6][4] * -32'h076) >> 8) + ((mcu[6][5] * -32'h0d0) >> 8) + ((mcu[6][6] * -32'h029) >> 8) + ((mcu[6][7] * 32'h0b0) >> 8) + ((mcu[7][0] * -32'h0d0) >> 8) + ((mcu[7][1] * 32'h030) >> 8) + ((mcu[7][2] * 32'h0f6) >> 8) + ((mcu[7][3] * 32'h08b) >> 8) + ((mcu[7][4] * -32'h08b) >> 8) + ((mcu[7][5] * -32'h0f6) >> 8) + ((mcu[7][6] * -32'h030) >> 8) + ((mcu[7][7] * 32'h0d0) >> 8);
	wire[63:0] cos14_term = ((mcu[0][0] * 32'h0b1) >> 8) + ((mcu[0][1] * -32'h0b1) >> 8) + ((mcu[0][2] * -32'h0b1) >> 8) + ((mcu[0][3] * 32'h0b1) >> 8) + ((mcu[0][4] * 32'h0b1) >> 8) + ((mcu[0][5] * -32'h0b1) >> 8) + ((mcu[0][6] * -32'h0b1) >> 8) + ((mcu[0][7] * 32'h0b1) >> 8) + ((mcu[1][0] * 32'h096) >> 8) + ((mcu[1][1] * -32'h096) >> 8) + ((mcu[1][2] * -32'h096) >> 8) + ((mcu[1][3] * 32'h096) >> 8) + ((mcu[1][4] * 32'h096) >> 8) + ((mcu[1][5] * -32'h096) >> 8) + ((mcu[1][6] * -32'h096) >> 8) + ((mcu[1][7] * 32'h096) >> 8) + ((mcu[2][0] * 32'h064) >> 8) + ((mcu[2][1] * -32'h064) >> 8) + ((mcu[2][2] * -32'h064) >> 8) + ((mcu[2][3] * 32'h064) >> 8) + ((mcu[2][4] * 32'h064) >> 8) + ((mcu[2][5] * -32'h064) >> 8) + ((mcu[2][6] * -32'h064) >> 8) + ((mcu[2][7] * 32'h064) >> 8) + ((mcu[3][0] * 32'h023) >> 8) + ((mcu[3][1] * -32'h023) >> 8) + ((mcu[3][2] * -32'h023) >> 8) + ((mcu[3][3] * 32'h023) >> 8) + ((mcu[3][4] * 32'h023) >> 8) + ((mcu[3][5] * -32'h023) >> 8) + ((mcu[3][6] * -32'h023) >> 8) + ((mcu[3][7] * 32'h023) >> 8) + ((mcu[4][0] * -32'h023) >> 8) + ((mcu[4][1] * 32'h023) >> 8) + ((mcu[4][2] * 32'h023) >> 8) + ((mcu[4][3] * -32'h023) >> 8) + ((mcu[4][4] * -32'h023) >> 8) + ((mcu[4][5] * 32'h023) >> 8) + ((mcu[4][6] * 32'h023) >> 8) + ((mcu[4][7] * -32'h023) >> 8) + ((mcu[5][0] * -32'h064) >> 8) + ((mcu[5][1] * 32'h064) >> 8) + ((mcu[5][2] * 32'h064) >> 8) + ((mcu[5][3] * -32'h064) >> 8) + ((mcu[5][4] * -32'h064) >> 8) + ((mcu[5][5] * 32'h064) >> 8) + ((mcu[5][6] * 32'h064) >> 8) + ((mcu[5][7] * -32'h064) >> 8) + ((mcu[6][0] * -32'h096) >> 8) + ((mcu[6][1] * 32'h096) >> 8) + ((mcu[6][2] * 32'h096) >> 8) + ((mcu[6][3] * -32'h096) >> 8) + ((mcu[6][4] * -32'h096) >> 8) + ((mcu[6][5] * 32'h096) >> 8) + ((mcu[6][6] * 32'h096) >> 8) + ((mcu[6][7] * -32'h096) >> 8) + ((mcu[7][0] * -32'h0b1) >> 8) + ((mcu[7][1] * 32'h0b1) >> 8) + ((mcu[7][2] * 32'h0b1) >> 8) + ((mcu[7][3] * -32'h0b1) >> 8) + ((mcu[7][4] * -32'h0b1) >> 8) + ((mcu[7][5] * 32'h0b1) >> 8) + ((mcu[7][6] * 32'h0b1) >> 8) + ((mcu[7][7] * -32'h0b1) >> 8);
	wire[63:0] cos15_term = ((mcu[0][0] * 32'h08b) >> 8) + ((mcu[0][1] * -32'h0f6) >> 8) + ((mcu[0][2] * 32'h030) >> 8) + ((mcu[0][3] * 32'h0d0) >> 8) + ((mcu[0][4] * -32'h0d0) >> 8) + ((mcu[0][5] * -32'h030) >> 8) + ((mcu[0][6] * 32'h0f6) >> 8) + ((mcu[0][7] * -32'h08b) >> 8) + ((mcu[1][0] * 32'h076) >> 8) + ((mcu[1][1] * -32'h0d0) >> 8) + ((mcu[1][2] * 32'h029) >> 8) + ((mcu[1][3] * 32'h0b0) >> 8) + ((mcu[1][4] * -32'h0b0) >> 8) + ((mcu[1][5] * -32'h029) >> 8) + ((mcu[1][6] * 32'h0d0) >> 8) + ((mcu[1][7] * -32'h076) >> 8) + ((mcu[2][0] * 32'h04f) >> 8) + ((mcu[2][1] * -32'h08b) >> 8) + ((mcu[2][2] * 32'h01b) >> 8) + ((mcu[2][3] * 32'h076) >> 8) + ((mcu[2][4] * -32'h076) >> 8) + ((mcu[2][5] * -32'h01b) >> 8) + ((mcu[2][6] * 32'h08b) >> 8) + ((mcu[2][7] * -32'h04f) >> 8) + ((mcu[3][0] * 32'h01b) >> 8) + ((mcu[3][1] * -32'h030) >> 8) + ((mcu[3][2] * 32'h009) >> 8) + ((mcu[3][3] * 32'h029) >> 8) + ((mcu[3][4] * -32'h029) >> 8) + ((mcu[3][5] * -32'h009) >> 8) + ((mcu[3][6] * 32'h030) >> 8) + ((mcu[3][7] * -32'h01b) >> 8) + ((mcu[4][0] * -32'h01b) >> 8) + ((mcu[4][1] * 32'h030) >> 8) + ((mcu[4][2] * -32'h009) >> 8) + ((mcu[4][3] * -32'h029) >> 8) + ((mcu[4][4] * 32'h029) >> 8) + ((mcu[4][5] * 32'h009) >> 8) + ((mcu[4][6] * -32'h030) >> 8) + ((mcu[4][7] * 32'h01b) >> 8) + ((mcu[5][0] * -32'h04f) >> 8) + ((mcu[5][1] * 32'h08b) >> 8) + ((mcu[5][2] * -32'h01b) >> 8) + ((mcu[5][3] * -32'h076) >> 8) + ((mcu[5][4] * 32'h076) >> 8) + ((mcu[5][5] * 32'h01b) >> 8) + ((mcu[5][6] * -32'h08b) >> 8) + ((mcu[5][7] * 32'h04f) >> 8) + ((mcu[6][0] * -32'h076) >> 8) + ((mcu[6][1] * 32'h0d0) >> 8) + ((mcu[6][2] * -32'h029) >> 8) + ((mcu[6][3] * -32'h0b0) >> 8) + ((mcu[6][4] * 32'h0b0) >> 8) + ((mcu[6][5] * 32'h029) >> 8) + ((mcu[6][6] * -32'h0d0) >> 8) + ((mcu[6][7] * 32'h076) >> 8) + ((mcu[7][0] * -32'h08b) >> 8) + ((mcu[7][1] * 32'h0f6) >> 8) + ((mcu[7][2] * -32'h030) >> 8) + ((mcu[7][3] * -32'h0d0) >> 8) + ((mcu[7][4] * 32'h0d0) >> 8) + ((mcu[7][5] * 32'h030) >> 8) + ((mcu[7][6] * -32'h0f6) >> 8) + ((mcu[7][7] * 32'h08b) >> 8);
	wire[63:0] cos16_term = ((mcu[0][0] * 32'h060) >> 8) + ((mcu[0][1] * -32'h0e7) >> 8) + ((mcu[0][2] * 32'h0e7) >> 8) + ((mcu[0][3] * -32'h060) >> 8) + ((mcu[0][4] * -32'h060) >> 8) + ((mcu[0][5] * 32'h0e7) >> 8) + ((mcu[0][6] * -32'h0e7) >> 8) + ((mcu[0][7] * 32'h060) >> 8) + ((mcu[1][0] * 32'h051) >> 8) + ((mcu[1][1] * -32'h0c4) >> 8) + ((mcu[1][2] * 32'h0c4) >> 8) + ((mcu[1][3] * -32'h051) >> 8) + ((mcu[1][4] * -32'h051) >> 8) + ((mcu[1][5] * 32'h0c4) >> 8) + ((mcu[1][6] * -32'h0c4) >> 8) + ((mcu[1][7] * 32'h051) >> 8) + ((mcu[2][0] * 32'h036) >> 8) + ((mcu[2][1] * -32'h083) >> 8) + ((mcu[2][2] * 32'h083) >> 8) + ((mcu[2][3] * -32'h036) >> 8) + ((mcu[2][4] * -32'h036) >> 8) + ((mcu[2][5] * 32'h083) >> 8) + ((mcu[2][6] * -32'h083) >> 8) + ((mcu[2][7] * 32'h036) >> 8) + ((mcu[3][0] * 32'h013) >> 8) + ((mcu[3][1] * -32'h02e) >> 8) + ((mcu[3][2] * 32'h02e) >> 8) + ((mcu[3][3] * -32'h013) >> 8) + ((mcu[3][4] * -32'h013) >> 8) + ((mcu[3][5] * 32'h02e) >> 8) + ((mcu[3][6] * -32'h02e) >> 8) + ((mcu[3][7] * 32'h013) >> 8) + ((mcu[4][0] * -32'h013) >> 8) + ((mcu[4][1] * 32'h02e) >> 8) + ((mcu[4][2] * -32'h02e) >> 8) + ((mcu[4][3] * 32'h013) >> 8) + ((mcu[4][4] * 32'h013) >> 8) + ((mcu[4][5] * -32'h02e) >> 8) + ((mcu[4][6] * 32'h02e) >> 8) + ((mcu[4][7] * -32'h013) >> 8) + ((mcu[5][0] * -32'h036) >> 8) + ((mcu[5][1] * 32'h083) >> 8) + ((mcu[5][2] * -32'h083) >> 8) + ((mcu[5][3] * 32'h036) >> 8) + ((mcu[5][4] * 32'h036) >> 8) + ((mcu[5][5] * -32'h083) >> 8) + ((mcu[5][6] * 32'h083) >> 8) + ((mcu[5][7] * -32'h036) >> 8) + ((mcu[6][0] * -32'h051) >> 8) + ((mcu[6][1] * 32'h0c4) >> 8) + ((mcu[6][2] * -32'h0c4) >> 8) + ((mcu[6][3] * 32'h051) >> 8) + ((mcu[6][4] * 32'h051) >> 8) + ((mcu[6][5] * -32'h0c4) >> 8) + ((mcu[6][6] * 32'h0c4) >> 8) + ((mcu[6][7] * -32'h051) >> 8) + ((mcu[7][0] * -32'h060) >> 8) + ((mcu[7][1] * 32'h0e7) >> 8) + ((mcu[7][2] * -32'h0e7) >> 8) + ((mcu[7][3] * 32'h060) >> 8) + ((mcu[7][4] * 32'h060) >> 8) + ((mcu[7][5] * -32'h0e7) >> 8) + ((mcu[7][6] * 32'h0e7) >> 8) + ((mcu[7][7] * -32'h060) >> 8);
	wire[63:0] cos17_term = ((mcu[0][0] * 32'h030) >> 8) + ((mcu[0][1] * -32'h08b) >> 8) + ((mcu[0][2] * 32'h0d0) >> 8) + ((mcu[0][3] * -32'h0f6) >> 8) + ((mcu[0][4] * 32'h0f6) >> 8) + ((mcu[0][5] * -32'h0d0) >> 8) + ((mcu[0][6] * 32'h08b) >> 8) + ((mcu[0][7] * -32'h030) >> 8) + ((mcu[1][0] * 32'h029) >> 8) + ((mcu[1][1] * -32'h076) >> 8) + ((mcu[1][2] * 32'h0b0) >> 8) + ((mcu[1][3] * -32'h0d0) >> 8) + ((mcu[1][4] * 32'h0d0) >> 8) + ((mcu[1][5] * -32'h0b0) >> 8) + ((mcu[1][6] * 32'h076) >> 8) + ((mcu[1][7] * -32'h029) >> 8) + ((mcu[2][0] * 32'h01b) >> 8) + ((mcu[2][1] * -32'h04f) >> 8) + ((mcu[2][2] * 32'h076) >> 8) + ((mcu[2][3] * -32'h08b) >> 8) + ((mcu[2][4] * 32'h08b) >> 8) + ((mcu[2][5] * -32'h076) >> 8) + ((mcu[2][6] * 32'h04f) >> 8) + ((mcu[2][7] * -32'h01b) >> 8) + ((mcu[3][0] * 32'h009) >> 8) + ((mcu[3][1] * -32'h01b) >> 8) + ((mcu[3][2] * 32'h029) >> 8) + ((mcu[3][3] * -32'h030) >> 8) + ((mcu[3][4] * 32'h030) >> 8) + ((mcu[3][5] * -32'h029) >> 8) + ((mcu[3][6] * 32'h01b) >> 8) + ((mcu[3][7] * -32'h009) >> 8) + ((mcu[4][0] * -32'h009) >> 8) + ((mcu[4][1] * 32'h01b) >> 8) + ((mcu[4][2] * -32'h029) >> 8) + ((mcu[4][3] * 32'h030) >> 8) + ((mcu[4][4] * -32'h030) >> 8) + ((mcu[4][5] * 32'h029) >> 8) + ((mcu[4][6] * -32'h01b) >> 8) + ((mcu[4][7] * 32'h009) >> 8) + ((mcu[5][0] * -32'h01b) >> 8) + ((mcu[5][1] * 32'h04f) >> 8) + ((mcu[5][2] * -32'h076) >> 8) + ((mcu[5][3] * 32'h08b) >> 8) + ((mcu[5][4] * -32'h08b) >> 8) + ((mcu[5][5] * 32'h076) >> 8) + ((mcu[5][6] * -32'h04f) >> 8) + ((mcu[5][7] * 32'h01b) >> 8) + ((mcu[6][0] * -32'h029) >> 8) + ((mcu[6][1] * 32'h076) >> 8) + ((mcu[6][2] * -32'h0b0) >> 8) + ((mcu[6][3] * 32'h0d0) >> 8) + ((mcu[6][4] * -32'h0d0) >> 8) + ((mcu[6][5] * 32'h0b0) >> 8) + ((mcu[6][6] * -32'h076) >> 8) + ((mcu[6][7] * 32'h029) >> 8) + ((mcu[7][0] * -32'h030) >> 8) + ((mcu[7][1] * 32'h08b) >> 8) + ((mcu[7][2] * -32'h0d0) >> 8) + ((mcu[7][3] * 32'h0f6) >> 8) + ((mcu[7][4] * -32'h0f6) >> 8) + ((mcu[7][5] * 32'h0d0) >> 8) + ((mcu[7][6] * -32'h08b) >> 8) + ((mcu[7][7] * 32'h030) >> 8);
	wire[63:0] cos20_term = ((mcu[0][0] * 32'h0ec) >> 8) + ((mcu[0][1] * 32'h0ec) >> 8) + ((mcu[0][2] * 32'h0ec) >> 8) + ((mcu[0][3] * 32'h0ec) >> 8) + ((mcu[0][4] * 32'h0ec) >> 8) + ((mcu[0][5] * 32'h0ec) >> 8) + ((mcu[0][6] * 32'h0ec) >> 8) + ((mcu[0][7] * 32'h0ec) >> 8) + ((mcu[1][0] * 32'h062) >> 8) + ((mcu[1][1] * 32'h062) >> 8) + ((mcu[1][2] * 32'h062) >> 8) + ((mcu[1][3] * 32'h062) >> 8) + ((mcu[1][4] * 32'h062) >> 8) + ((mcu[1][5] * 32'h062) >> 8) + ((mcu[1][6] * 32'h062) >> 8) + ((mcu[1][7] * 32'h062) >> 8) + ((mcu[2][0] * -32'h062) >> 8) + ((mcu[2][1] * -32'h062) >> 8) + ((mcu[2][2] * -32'h062) >> 8) + ((mcu[2][3] * -32'h062) >> 8) + ((mcu[2][4] * -32'h062) >> 8) + ((mcu[2][5] * -32'h062) >> 8) + ((mcu[2][6] * -32'h062) >> 8) + ((mcu[2][7] * -32'h062) >> 8) + ((mcu[3][0] * -32'h0ec) >> 8) + ((mcu[3][1] * -32'h0ec) >> 8) + ((mcu[3][2] * -32'h0ec) >> 8) + ((mcu[3][3] * -32'h0ec) >> 8) + ((mcu[3][4] * -32'h0ec) >> 8) + ((mcu[3][5] * -32'h0ec) >> 8) + ((mcu[3][6] * -32'h0ec) >> 8) + ((mcu[3][7] * -32'h0ec) >> 8) + ((mcu[4][0] * -32'h0ec) >> 8) + ((mcu[4][1] * -32'h0ec) >> 8) + ((mcu[4][2] * -32'h0ec) >> 8) + ((mcu[4][3] * -32'h0ec) >> 8) + ((mcu[4][4] * -32'h0ec) >> 8) + ((mcu[4][5] * -32'h0ec) >> 8) + ((mcu[4][6] * -32'h0ec) >> 8) + ((mcu[4][7] * -32'h0ec) >> 8) + ((mcu[5][0] * -32'h062) >> 8) + ((mcu[5][1] * -32'h062) >> 8) + ((mcu[5][2] * -32'h062) >> 8) + ((mcu[5][3] * -32'h062) >> 8) + ((mcu[5][4] * -32'h062) >> 8) + ((mcu[5][5] * -32'h062) >> 8) + ((mcu[5][6] * -32'h062) >> 8) + ((mcu[5][7] * -32'h062) >> 8) + ((mcu[6][0] * 32'h062) >> 8) + ((mcu[6][1] * 32'h062) >> 8) + ((mcu[6][2] * 32'h062) >> 8) + ((mcu[6][3] * 32'h062) >> 8) + ((mcu[6][4] * 32'h062) >> 8) + ((mcu[6][5] * 32'h062) >> 8) + ((mcu[6][6] * 32'h062) >> 8) + ((mcu[6][7] * 32'h062) >> 8) + ((mcu[7][0] * 32'h0ec) >> 8) + ((mcu[7][1] * 32'h0ec) >> 8) + ((mcu[7][2] * 32'h0ec) >> 8) + ((mcu[7][3] * 32'h0ec) >> 8) + ((mcu[7][4] * 32'h0ec) >> 8) + ((mcu[7][5] * 32'h0ec) >> 8) + ((mcu[7][6] * 32'h0ec) >> 8) + ((mcu[7][7] * 32'h0ec) >> 8);
	wire[63:0] cos21_term = ((mcu[0][0] * 32'h0e7) >> 8) + ((mcu[0][1] * 32'h0c4) >> 8) + ((mcu[0][2] * 32'h083) >> 8) + ((mcu[0][3] * 32'h02e) >> 8) + ((mcu[0][4] * -32'h02e) >> 8) + ((mcu[0][5] * -32'h083) >> 8) + ((mcu[0][6] * -32'h0c4) >> 8) + ((mcu[0][7] * -32'h0e7) >> 8) + ((mcu[1][0] * 32'h060) >> 8) + ((mcu[1][1] * 32'h051) >> 8) + ((mcu[1][2] * 32'h036) >> 8) + ((mcu[1][3] * 32'h013) >> 8) + ((mcu[1][4] * -32'h013) >> 8) + ((mcu[1][5] * -32'h036) >> 8) + ((mcu[1][6] * -32'h051) >> 8) + ((mcu[1][7] * -32'h060) >> 8) + ((mcu[2][0] * -32'h060) >> 8) + ((mcu[2][1] * -32'h051) >> 8) + ((mcu[2][2] * -32'h036) >> 8) + ((mcu[2][3] * -32'h013) >> 8) + ((mcu[2][4] * 32'h013) >> 8) + ((mcu[2][5] * 32'h036) >> 8) + ((mcu[2][6] * 32'h051) >> 8) + ((mcu[2][7] * 32'h060) >> 8) + ((mcu[3][0] * -32'h0e7) >> 8) + ((mcu[3][1] * -32'h0c4) >> 8) + ((mcu[3][2] * -32'h083) >> 8) + ((mcu[3][3] * -32'h02e) >> 8) + ((mcu[3][4] * 32'h02e) >> 8) + ((mcu[3][5] * 32'h083) >> 8) + ((mcu[3][6] * 32'h0c4) >> 8) + ((mcu[3][7] * 32'h0e7) >> 8) + ((mcu[4][0] * -32'h0e7) >> 8) + ((mcu[4][1] * -32'h0c4) >> 8) + ((mcu[4][2] * -32'h083) >> 8) + ((mcu[4][3] * -32'h02e) >> 8) + ((mcu[4][4] * 32'h02e) >> 8) + ((mcu[4][5] * 32'h083) >> 8) + ((mcu[4][6] * 32'h0c4) >> 8) + ((mcu[4][7] * 32'h0e7) >> 8) + ((mcu[5][0] * -32'h060) >> 8) + ((mcu[5][1] * -32'h051) >> 8) + ((mcu[5][2] * -32'h036) >> 8) + ((mcu[5][3] * -32'h013) >> 8) + ((mcu[5][4] * 32'h013) >> 8) + ((mcu[5][5] * 32'h036) >> 8) + ((mcu[5][6] * 32'h051) >> 8) + ((mcu[5][7] * 32'h060) >> 8) + ((mcu[6][0] * 32'h060) >> 8) + ((mcu[6][1] * 32'h051) >> 8) + ((mcu[6][2] * 32'h036) >> 8) + ((mcu[6][3] * 32'h013) >> 8) + ((mcu[6][4] * -32'h013) >> 8) + ((mcu[6][5] * -32'h036) >> 8) + ((mcu[6][6] * -32'h051) >> 8) + ((mcu[6][7] * -32'h060) >> 8) + ((mcu[7][0] * 32'h0e7) >> 8) + ((mcu[7][1] * 32'h0c4) >> 8) + ((mcu[7][2] * 32'h083) >> 8) + ((mcu[7][3] * 32'h02e) >> 8) + ((mcu[7][4] * -32'h02e) >> 8) + ((mcu[7][5] * -32'h083) >> 8) + ((mcu[7][6] * -32'h0c4) >> 8) + ((mcu[7][7] * -32'h0e7) >> 8);
	wire[63:0] cos22_term = ((mcu[0][0] * 32'h0da) >> 8) + ((mcu[0][1] * 32'h05a) >> 8) + ((mcu[0][2] * -32'h05a) >> 8) + ((mcu[0][3] * -32'h0da) >> 8) + ((mcu[0][4] * -32'h0da) >> 8) + ((mcu[0][5] * -32'h05a) >> 8) + ((mcu[0][6] * 32'h05a) >> 8) + ((mcu[0][7] * 32'h0da) >> 8) + ((mcu[1][0] * 32'h05a) >> 8) + ((mcu[1][1] * 32'h025) >> 8) + ((mcu[1][2] * -32'h025) >> 8) + ((mcu[1][3] * -32'h05a) >> 8) + ((mcu[1][4] * -32'h05a) >> 8) + ((mcu[1][5] * -32'h025) >> 8) + ((mcu[1][6] * 32'h025) >> 8) + ((mcu[1][7] * 32'h05a) >> 8) + ((mcu[2][0] * -32'h05a) >> 8) + ((mcu[2][1] * -32'h025) >> 8) + ((mcu[2][2] * 32'h025) >> 8) + ((mcu[2][3] * 32'h05a) >> 8) + ((mcu[2][4] * 32'h05a) >> 8) + ((mcu[2][5] * 32'h025) >> 8) + ((mcu[2][6] * -32'h025) >> 8) + ((mcu[2][7] * -32'h05a) >> 8) + ((mcu[3][0] * -32'h0da) >> 8) + ((mcu[3][1] * -32'h05a) >> 8) + ((mcu[3][2] * 32'h05a) >> 8) + ((mcu[3][3] * 32'h0da) >> 8) + ((mcu[3][4] * 32'h0da) >> 8) + ((mcu[3][5] * 32'h05a) >> 8) + ((mcu[3][6] * -32'h05a) >> 8) + ((mcu[3][7] * -32'h0da) >> 8) + ((mcu[4][0] * -32'h0da) >> 8) + ((mcu[4][1] * -32'h05a) >> 8) + ((mcu[4][2] * 32'h05a) >> 8) + ((mcu[4][3] * 32'h0da) >> 8) + ((mcu[4][4] * 32'h0da) >> 8) + ((mcu[4][5] * 32'h05a) >> 8) + ((mcu[4][6] * -32'h05a) >> 8) + ((mcu[4][7] * -32'h0da) >> 8) + ((mcu[5][0] * -32'h05a) >> 8) + ((mcu[5][1] * -32'h025) >> 8) + ((mcu[5][2] * 32'h025) >> 8) + ((mcu[5][3] * 32'h05a) >> 8) + ((mcu[5][4] * 32'h05a) >> 8) + ((mcu[5][5] * 32'h025) >> 8) + ((mcu[5][6] * -32'h025) >> 8) + ((mcu[5][7] * -32'h05a) >> 8) + ((mcu[6][0] * 32'h05a) >> 8) + ((mcu[6][1] * 32'h025) >> 8) + ((mcu[6][2] * -32'h025) >> 8) + ((mcu[6][3] * -32'h05a) >> 8) + ((mcu[6][4] * -32'h05a) >> 8) + ((mcu[6][5] * -32'h025) >> 8) + ((mcu[6][6] * 32'h025) >> 8) + ((mcu[6][7] * 32'h05a) >> 8) + ((mcu[7][0] * 32'h0da) >> 8) + ((mcu[7][1] * 32'h05a) >> 8) + ((mcu[7][2] * -32'h05a) >> 8) + ((mcu[7][3] * -32'h0da) >> 8) + ((mcu[7][4] * -32'h0da) >> 8) + ((mcu[7][5] * -32'h05a) >> 8) + ((mcu[7][6] * 32'h05a) >> 8) + ((mcu[7][7] * 32'h0da) >> 8);
	wire[63:0] cos23_term = ((mcu[0][0] * 32'h0c4) >> 8) + ((mcu[0][1] * -32'h02e) >> 8) + ((mcu[0][2] * -32'h0e7) >> 8) + ((mcu[0][3] * -32'h083) >> 8) + ((mcu[0][4] * 32'h083) >> 8) + ((mcu[0][5] * 32'h0e7) >> 8) + ((mcu[0][6] * 32'h02e) >> 8) + ((mcu[0][7] * -32'h0c4) >> 8) + ((mcu[1][0] * 32'h051) >> 8) + ((mcu[1][1] * -32'h013) >> 8) + ((mcu[1][2] * -32'h060) >> 8) + ((mcu[1][3] * -32'h036) >> 8) + ((mcu[1][4] * 32'h036) >> 8) + ((mcu[1][5] * 32'h060) >> 8) + ((mcu[1][6] * 32'h013) >> 8) + ((mcu[1][7] * -32'h051) >> 8) + ((mcu[2][0] * -32'h051) >> 8) + ((mcu[2][1] * 32'h013) >> 8) + ((mcu[2][2] * 32'h060) >> 8) + ((mcu[2][3] * 32'h036) >> 8) + ((mcu[2][4] * -32'h036) >> 8) + ((mcu[2][5] * -32'h060) >> 8) + ((mcu[2][6] * -32'h013) >> 8) + ((mcu[2][7] * 32'h051) >> 8) + ((mcu[3][0] * -32'h0c4) >> 8) + ((mcu[3][1] * 32'h02e) >> 8) + ((mcu[3][2] * 32'h0e7) >> 8) + ((mcu[3][3] * 32'h083) >> 8) + ((mcu[3][4] * -32'h083) >> 8) + ((mcu[3][5] * -32'h0e7) >> 8) + ((mcu[3][6] * -32'h02e) >> 8) + ((mcu[3][7] * 32'h0c4) >> 8) + ((mcu[4][0] * -32'h0c4) >> 8) + ((mcu[4][1] * 32'h02e) >> 8) + ((mcu[4][2] * 32'h0e7) >> 8) + ((mcu[4][3] * 32'h083) >> 8) + ((mcu[4][4] * -32'h083) >> 8) + ((mcu[4][5] * -32'h0e7) >> 8) + ((mcu[4][6] * -32'h02e) >> 8) + ((mcu[4][7] * 32'h0c4) >> 8) + ((mcu[5][0] * -32'h051) >> 8) + ((mcu[5][1] * 32'h013) >> 8) + ((mcu[5][2] * 32'h060) >> 8) + ((mcu[5][3] * 32'h036) >> 8) + ((mcu[5][4] * -32'h036) >> 8) + ((mcu[5][5] * -32'h060) >> 8) + ((mcu[5][6] * -32'h013) >> 8) + ((mcu[5][7] * 32'h051) >> 8) + ((mcu[6][0] * 32'h051) >> 8) + ((mcu[6][1] * -32'h013) >> 8) + ((mcu[6][2] * -32'h060) >> 8) + ((mcu[6][3] * -32'h036) >> 8) + ((mcu[6][4] * 32'h036) >> 8) + ((mcu[6][5] * 32'h060) >> 8) + ((mcu[6][6] * 32'h013) >> 8) + ((mcu[6][7] * -32'h051) >> 8) + ((mcu[7][0] * 32'h0c4) >> 8) + ((mcu[7][1] * -32'h02e) >> 8) + ((mcu[7][2] * -32'h0e7) >> 8) + ((mcu[7][3] * -32'h083) >> 8) + ((mcu[7][4] * 32'h083) >> 8) + ((mcu[7][5] * 32'h0e7) >> 8) + ((mcu[7][6] * 32'h02e) >> 8) + ((mcu[7][7] * -32'h0c4) >> 8);
	wire[63:0] cos24_term = ((mcu[0][0] * 32'h0a7) >> 8) + ((mcu[0][1] * -32'h0a7) >> 8) + ((mcu[0][2] * -32'h0a7) >> 8) + ((mcu[0][3] * 32'h0a7) >> 8) + ((mcu[0][4] * 32'h0a7) >> 8) + ((mcu[0][5] * -32'h0a7) >> 8) + ((mcu[0][6] * -32'h0a7) >> 8) + ((mcu[0][7] * 32'h0a7) >> 8) + ((mcu[1][0] * 32'h045) >> 8) + ((mcu[1][1] * -32'h045) >> 8) + ((mcu[1][2] * -32'h045) >> 8) + ((mcu[1][3] * 32'h045) >> 8) + ((mcu[1][4] * 32'h045) >> 8) + ((mcu[1][5] * -32'h045) >> 8) + ((mcu[1][6] * -32'h045) >> 8) + ((mcu[1][7] * 32'h045) >> 8) + ((mcu[2][0] * -32'h045) >> 8) + ((mcu[2][1] * 32'h045) >> 8) + ((mcu[2][2] * 32'h045) >> 8) + ((mcu[2][3] * -32'h045) >> 8) + ((mcu[2][4] * -32'h045) >> 8) + ((mcu[2][5] * 32'h045) >> 8) + ((mcu[2][6] * 32'h045) >> 8) + ((mcu[2][7] * -32'h045) >> 8) + ((mcu[3][0] * -32'h0a7) >> 8) + ((mcu[3][1] * 32'h0a7) >> 8) + ((mcu[3][2] * 32'h0a7) >> 8) + ((mcu[3][3] * -32'h0a7) >> 8) + ((mcu[3][4] * -32'h0a7) >> 8) + ((mcu[3][5] * 32'h0a7) >> 8) + ((mcu[3][6] * 32'h0a7) >> 8) + ((mcu[3][7] * -32'h0a7) >> 8) + ((mcu[4][0] * -32'h0a7) >> 8) + ((mcu[4][1] * 32'h0a7) >> 8) + ((mcu[4][2] * 32'h0a7) >> 8) + ((mcu[4][3] * -32'h0a7) >> 8) + ((mcu[4][4] * -32'h0a7) >> 8) + ((mcu[4][5] * 32'h0a7) >> 8) + ((mcu[4][6] * 32'h0a7) >> 8) + ((mcu[4][7] * -32'h0a7) >> 8) + ((mcu[5][0] * -32'h045) >> 8) + ((mcu[5][1] * 32'h045) >> 8) + ((mcu[5][2] * 32'h045) >> 8) + ((mcu[5][3] * -32'h045) >> 8) + ((mcu[5][4] * -32'h045) >> 8) + ((mcu[5][5] * 32'h045) >> 8) + ((mcu[5][6] * 32'h045) >> 8) + ((mcu[5][7] * -32'h045) >> 8) + ((mcu[6][0] * 32'h045) >> 8) + ((mcu[6][1] * -32'h045) >> 8) + ((mcu[6][2] * -32'h045) >> 8) + ((mcu[6][3] * 32'h045) >> 8) + ((mcu[6][4] * 32'h045) >> 8) + ((mcu[6][5] * -32'h045) >> 8) + ((mcu[6][6] * -32'h045) >> 8) + ((mcu[6][7] * 32'h045) >> 8) + ((mcu[7][0] * 32'h0a7) >> 8) + ((mcu[7][1] * -32'h0a7) >> 8) + ((mcu[7][2] * -32'h0a7) >> 8) + ((mcu[7][3] * 32'h0a7) >> 8) + ((mcu[7][4] * 32'h0a7) >> 8) + ((mcu[7][5] * -32'h0a7) >> 8) + ((mcu[7][6] * -32'h0a7) >> 8) + ((mcu[7][7] * 32'h0a7) >> 8);
	wire[63:0] cos25_term = ((mcu[0][0] * 32'h083) >> 8) + ((mcu[0][1] * -32'h0e7) >> 8) + ((mcu[0][2] * 32'h02e) >> 8) + ((mcu[0][3] * 32'h0c4) >> 8) + ((mcu[0][4] * -32'h0c4) >> 8) + ((mcu[0][5] * -32'h02e) >> 8) + ((mcu[0][6] * 32'h0e7) >> 8) + ((mcu[0][7] * -32'h083) >> 8) + ((mcu[1][0] * 32'h036) >> 8) + ((mcu[1][1] * -32'h060) >> 8) + ((mcu[1][2] * 32'h013) >> 8) + ((mcu[1][3] * 32'h051) >> 8) + ((mcu[1][4] * -32'h051) >> 8) + ((mcu[1][5] * -32'h013) >> 8) + ((mcu[1][6] * 32'h060) >> 8) + ((mcu[1][7] * -32'h036) >> 8) + ((mcu[2][0] * -32'h036) >> 8) + ((mcu[2][1] * 32'h060) >> 8) + ((mcu[2][2] * -32'h013) >> 8) + ((mcu[2][3] * -32'h051) >> 8) + ((mcu[2][4] * 32'h051) >> 8) + ((mcu[2][5] * 32'h013) >> 8) + ((mcu[2][6] * -32'h060) >> 8) + ((mcu[2][7] * 32'h036) >> 8) + ((mcu[3][0] * -32'h083) >> 8) + ((mcu[3][1] * 32'h0e7) >> 8) + ((mcu[3][2] * -32'h02e) >> 8) + ((mcu[3][3] * -32'h0c4) >> 8) + ((mcu[3][4] * 32'h0c4) >> 8) + ((mcu[3][5] * 32'h02e) >> 8) + ((mcu[3][6] * -32'h0e7) >> 8) + ((mcu[3][7] * 32'h083) >> 8) + ((mcu[4][0] * -32'h083) >> 8) + ((mcu[4][1] * 32'h0e7) >> 8) + ((mcu[4][2] * -32'h02e) >> 8) + ((mcu[4][3] * -32'h0c4) >> 8) + ((mcu[4][4] * 32'h0c4) >> 8) + ((mcu[4][5] * 32'h02e) >> 8) + ((mcu[4][6] * -32'h0e7) >> 8) + ((mcu[4][7] * 32'h083) >> 8) + ((mcu[5][0] * -32'h036) >> 8) + ((mcu[5][1] * 32'h060) >> 8) + ((mcu[5][2] * -32'h013) >> 8) + ((mcu[5][3] * -32'h051) >> 8) + ((mcu[5][4] * 32'h051) >> 8) + ((mcu[5][5] * 32'h013) >> 8) + ((mcu[5][6] * -32'h060) >> 8) + ((mcu[5][7] * 32'h036) >> 8) + ((mcu[6][0] * 32'h036) >> 8) + ((mcu[6][1] * -32'h060) >> 8) + ((mcu[6][2] * 32'h013) >> 8) + ((mcu[6][3] * 32'h051) >> 8) + ((mcu[6][4] * -32'h051) >> 8) + ((mcu[6][5] * -32'h013) >> 8) + ((mcu[6][6] * 32'h060) >> 8) + ((mcu[6][7] * -32'h036) >> 8) + ((mcu[7][0] * 32'h083) >> 8) + ((mcu[7][1] * -32'h0e7) >> 8) + ((mcu[7][2] * 32'h02e) >> 8) + ((mcu[7][3] * 32'h0c4) >> 8) + ((mcu[7][4] * -32'h0c4) >> 8) + ((mcu[7][5] * -32'h02e) >> 8) + ((mcu[7][6] * 32'h0e7) >> 8) + ((mcu[7][7] * -32'h083) >> 8);
	wire[63:0] cos26_term = ((mcu[0][0] * 32'h05a) >> 8) + ((mcu[0][1] * -32'h0da) >> 8) + ((mcu[0][2] * 32'h0da) >> 8) + ((mcu[0][3] * -32'h05a) >> 8) + ((mcu[0][4] * -32'h05a) >> 8) + ((mcu[0][5] * 32'h0da) >> 8) + ((mcu[0][6] * -32'h0da) >> 8) + ((mcu[0][7] * 32'h05a) >> 8) + ((mcu[1][0] * 32'h025) >> 8) + ((mcu[1][1] * -32'h05a) >> 8) + ((mcu[1][2] * 32'h05a) >> 8) + ((mcu[1][3] * -32'h025) >> 8) + ((mcu[1][4] * -32'h025) >> 8) + ((mcu[1][5] * 32'h05a) >> 8) + ((mcu[1][6] * -32'h05a) >> 8) + ((mcu[1][7] * 32'h025) >> 8) + ((mcu[2][0] * -32'h025) >> 8) + ((mcu[2][1] * 32'h05a) >> 8) + ((mcu[2][2] * -32'h05a) >> 8) + ((mcu[2][3] * 32'h025) >> 8) + ((mcu[2][4] * 32'h025) >> 8) + ((mcu[2][5] * -32'h05a) >> 8) + ((mcu[2][6] * 32'h05a) >> 8) + ((mcu[2][7] * -32'h025) >> 8) + ((mcu[3][0] * -32'h05a) >> 8) + ((mcu[3][1] * 32'h0da) >> 8) + ((mcu[3][2] * -32'h0da) >> 8) + ((mcu[3][3] * 32'h05a) >> 8) + ((mcu[3][4] * 32'h05a) >> 8) + ((mcu[3][5] * -32'h0da) >> 8) + ((mcu[3][6] * 32'h0da) >> 8) + ((mcu[3][7] * -32'h05a) >> 8) + ((mcu[4][0] * -32'h05a) >> 8) + ((mcu[4][1] * 32'h0da) >> 8) + ((mcu[4][2] * -32'h0da) >> 8) + ((mcu[4][3] * 32'h05a) >> 8) + ((mcu[4][4] * 32'h05a) >> 8) + ((mcu[4][5] * -32'h0da) >> 8) + ((mcu[4][6] * 32'h0da) >> 8) + ((mcu[4][7] * -32'h05a) >> 8) + ((mcu[5][0] * -32'h025) >> 8) + ((mcu[5][1] * 32'h05a) >> 8) + ((mcu[5][2] * -32'h05a) >> 8) + ((mcu[5][3] * 32'h025) >> 8) + ((mcu[5][4] * 32'h025) >> 8) + ((mcu[5][5] * -32'h05a) >> 8) + ((mcu[5][6] * 32'h05a) >> 8) + ((mcu[5][7] * -32'h025) >> 8) + ((mcu[6][0] * 32'h025) >> 8) + ((mcu[6][1] * -32'h05a) >> 8) + ((mcu[6][2] * 32'h05a) >> 8) + ((mcu[6][3] * -32'h025) >> 8) + ((mcu[6][4] * -32'h025) >> 8) + ((mcu[6][5] * 32'h05a) >> 8) + ((mcu[6][6] * -32'h05a) >> 8) + ((mcu[6][7] * 32'h025) >> 8) + ((mcu[7][0] * 32'h05a) >> 8) + ((mcu[7][1] * -32'h0da) >> 8) + ((mcu[7][2] * 32'h0da) >> 8) + ((mcu[7][3] * -32'h05a) >> 8) + ((mcu[7][4] * -32'h05a) >> 8) + ((mcu[7][5] * 32'h0da) >> 8) + ((mcu[7][6] * -32'h0da) >> 8) + ((mcu[7][7] * 32'h05a) >> 8);
	wire[63:0] cos27_term = ((mcu[0][0] * 32'h02e) >> 8) + ((mcu[0][1] * -32'h083) >> 8) + ((mcu[0][2] * 32'h0c4) >> 8) + ((mcu[0][3] * -32'h0e7) >> 8) + ((mcu[0][4] * 32'h0e7) >> 8) + ((mcu[0][5] * -32'h0c4) >> 8) + ((mcu[0][6] * 32'h083) >> 8) + ((mcu[0][7] * -32'h02e) >> 8) + ((mcu[1][0] * 32'h013) >> 8) + ((mcu[1][1] * -32'h036) >> 8) + ((mcu[1][2] * 32'h051) >> 8) + ((mcu[1][3] * -32'h060) >> 8) + ((mcu[1][4] * 32'h060) >> 8) + ((mcu[1][5] * -32'h051) >> 8) + ((mcu[1][6] * 32'h036) >> 8) + ((mcu[1][7] * -32'h013) >> 8) + ((mcu[2][0] * -32'h013) >> 8) + ((mcu[2][1] * 32'h036) >> 8) + ((mcu[2][2] * -32'h051) >> 8) + ((mcu[2][3] * 32'h060) >> 8) + ((mcu[2][4] * -32'h060) >> 8) + ((mcu[2][5] * 32'h051) >> 8) + ((mcu[2][6] * -32'h036) >> 8) + ((mcu[2][7] * 32'h013) >> 8) + ((mcu[3][0] * -32'h02e) >> 8) + ((mcu[3][1] * 32'h083) >> 8) + ((mcu[3][2] * -32'h0c4) >> 8) + ((mcu[3][3] * 32'h0e7) >> 8) + ((mcu[3][4] * -32'h0e7) >> 8) + ((mcu[3][5] * 32'h0c4) >> 8) + ((mcu[3][6] * -32'h083) >> 8) + ((mcu[3][7] * 32'h02e) >> 8) + ((mcu[4][0] * -32'h02e) >> 8) + ((mcu[4][1] * 32'h083) >> 8) + ((mcu[4][2] * -32'h0c4) >> 8) + ((mcu[4][3] * 32'h0e7) >> 8) + ((mcu[4][4] * -32'h0e7) >> 8) + ((mcu[4][5] * 32'h0c4) >> 8) + ((mcu[4][6] * -32'h083) >> 8) + ((mcu[4][7] * 32'h02e) >> 8) + ((mcu[5][0] * -32'h013) >> 8) + ((mcu[5][1] * 32'h036) >> 8) + ((mcu[5][2] * -32'h051) >> 8) + ((mcu[5][3] * 32'h060) >> 8) + ((mcu[5][4] * -32'h060) >> 8) + ((mcu[5][5] * 32'h051) >> 8) + ((mcu[5][6] * -32'h036) >> 8) + ((mcu[5][7] * 32'h013) >> 8) + ((mcu[6][0] * 32'h013) >> 8) + ((mcu[6][1] * -32'h036) >> 8) + ((mcu[6][2] * 32'h051) >> 8) + ((mcu[6][3] * -32'h060) >> 8) + ((mcu[6][4] * 32'h060) >> 8) + ((mcu[6][5] * -32'h051) >> 8) + ((mcu[6][6] * 32'h036) >> 8) + ((mcu[6][7] * -32'h013) >> 8) + ((mcu[7][0] * 32'h02e) >> 8) + ((mcu[7][1] * -32'h083) >> 8) + ((mcu[7][2] * 32'h0c4) >> 8) + ((mcu[7][3] * -32'h0e7) >> 8) + ((mcu[7][4] * 32'h0e7) >> 8) + ((mcu[7][5] * -32'h0c4) >> 8) + ((mcu[7][6] * 32'h083) >> 8) + ((mcu[7][7] * -32'h02e) >> 8);
	wire[63:0] cos30_term = ((mcu[0][0] * 32'h0d4) >> 8) + ((mcu[0][1] * 32'h0d4) >> 8) + ((mcu[0][2] * 32'h0d4) >> 8) + ((mcu[0][3] * 32'h0d4) >> 8) + ((mcu[0][4] * 32'h0d4) >> 8) + ((mcu[0][5] * 32'h0d4) >> 8) + ((mcu[0][6] * 32'h0d4) >> 8) + ((mcu[0][7] * 32'h0d4) >> 8) + ((mcu[1][0] * -32'h031) >> 8) + ((mcu[1][1] * -32'h031) >> 8) + ((mcu[1][2] * -32'h031) >> 8) + ((mcu[1][3] * -32'h031) >> 8) + ((mcu[1][4] * -32'h031) >> 8) + ((mcu[1][5] * -32'h031) >> 8) + ((mcu[1][6] * -32'h031) >> 8) + ((mcu[1][7] * -32'h031) >> 8) + ((mcu[2][0] * -32'h0fb) >> 8) + ((mcu[2][1] * -32'h0fb) >> 8) + ((mcu[2][2] * -32'h0fb) >> 8) + ((mcu[2][3] * -32'h0fb) >> 8) + ((mcu[2][4] * -32'h0fb) >> 8) + ((mcu[2][5] * -32'h0fb) >> 8) + ((mcu[2][6] * -32'h0fb) >> 8) + ((mcu[2][7] * -32'h0fb) >> 8) + ((mcu[3][0] * -32'h08e) >> 8) + ((mcu[3][1] * -32'h08e) >> 8) + ((mcu[3][2] * -32'h08e) >> 8) + ((mcu[3][3] * -32'h08e) >> 8) + ((mcu[3][4] * -32'h08e) >> 8) + ((mcu[3][5] * -32'h08e) >> 8) + ((mcu[3][6] * -32'h08e) >> 8) + ((mcu[3][7] * -32'h08e) >> 8) + ((mcu[4][0] * 32'h08e) >> 8) + ((mcu[4][1] * 32'h08e) >> 8) + ((mcu[4][2] * 32'h08e) >> 8) + ((mcu[4][3] * 32'h08e) >> 8) + ((mcu[4][4] * 32'h08e) >> 8) + ((mcu[4][5] * 32'h08e) >> 8) + ((mcu[4][6] * 32'h08e) >> 8) + ((mcu[4][7] * 32'h08e) >> 8) + ((mcu[5][0] * 32'h0fb) >> 8) + ((mcu[5][1] * 32'h0fb) >> 8) + ((mcu[5][2] * 32'h0fb) >> 8) + ((mcu[5][3] * 32'h0fb) >> 8) + ((mcu[5][4] * 32'h0fb) >> 8) + ((mcu[5][5] * 32'h0fb) >> 8) + ((mcu[5][6] * 32'h0fb) >> 8) + ((mcu[5][7] * 32'h0fb) >> 8) + ((mcu[6][0] * 32'h031) >> 8) + ((mcu[6][1] * 32'h031) >> 8) + ((mcu[6][2] * 32'h031) >> 8) + ((mcu[6][3] * 32'h031) >> 8) + ((mcu[6][4] * 32'h031) >> 8) + ((mcu[6][5] * 32'h031) >> 8) + ((mcu[6][6] * 32'h031) >> 8) + ((mcu[6][7] * 32'h031) >> 8) + ((mcu[7][0] * -32'h0d4) >> 8) + ((mcu[7][1] * -32'h0d4) >> 8) + ((mcu[7][2] * -32'h0d4) >> 8) + ((mcu[7][3] * -32'h0d4) >> 8) + ((mcu[7][4] * -32'h0d4) >> 8) + ((mcu[7][5] * -32'h0d4) >> 8) + ((mcu[7][6] * -32'h0d4) >> 8) + ((mcu[7][7] * -32'h0d4) >> 8);
	wire[63:0] cos31_term = ((mcu[0][0] * 32'h0d0) >> 8) + ((mcu[0][1] * 32'h0b0) >> 8) + ((mcu[0][2] * 32'h076) >> 8) + ((mcu[0][3] * 32'h029) >> 8) + ((mcu[0][4] * -32'h029) >> 8) + ((mcu[0][5] * -32'h076) >> 8) + ((mcu[0][6] * -32'h0b0) >> 8) + ((mcu[0][7] * -32'h0d0) >> 8) + ((mcu[1][0] * -32'h030) >> 8) + ((mcu[1][1] * -32'h029) >> 8) + ((mcu[1][2] * -32'h01b) >> 8) + ((mcu[1][3] * -32'h009) >> 8) + ((mcu[1][4] * 32'h009) >> 8) + ((mcu[1][5] * 32'h01b) >> 8) + ((mcu[1][6] * 32'h029) >> 8) + ((mcu[1][7] * 32'h030) >> 8) + ((mcu[2][0] * -32'h0f6) >> 8) + ((mcu[2][1] * -32'h0d0) >> 8) + ((mcu[2][2] * -32'h08b) >> 8) + ((mcu[2][3] * -32'h030) >> 8) + ((mcu[2][4] * 32'h030) >> 8) + ((mcu[2][5] * 32'h08b) >> 8) + ((mcu[2][6] * 32'h0d0) >> 8) + ((mcu[2][7] * 32'h0f6) >> 8) + ((mcu[3][0] * -32'h08b) >> 8) + ((mcu[3][1] * -32'h076) >> 8) + ((mcu[3][2] * -32'h04f) >> 8) + ((mcu[3][3] * -32'h01b) >> 8) + ((mcu[3][4] * 32'h01b) >> 8) + ((mcu[3][5] * 32'h04f) >> 8) + ((mcu[3][6] * 32'h076) >> 8) + ((mcu[3][7] * 32'h08b) >> 8) + ((mcu[4][0] * 32'h08b) >> 8) + ((mcu[4][1] * 32'h076) >> 8) + ((mcu[4][2] * 32'h04f) >> 8) + ((mcu[4][3] * 32'h01b) >> 8) + ((mcu[4][4] * -32'h01b) >> 8) + ((mcu[4][5] * -32'h04f) >> 8) + ((mcu[4][6] * -32'h076) >> 8) + ((mcu[4][7] * -32'h08b) >> 8) + ((mcu[5][0] * 32'h0f6) >> 8) + ((mcu[5][1] * 32'h0d0) >> 8) + ((mcu[5][2] * 32'h08b) >> 8) + ((mcu[5][3] * 32'h030) >> 8) + ((mcu[5][4] * -32'h030) >> 8) + ((mcu[5][5] * -32'h08b) >> 8) + ((mcu[5][6] * -32'h0d0) >> 8) + ((mcu[5][7] * -32'h0f6) >> 8) + ((mcu[6][0] * 32'h030) >> 8) + ((mcu[6][1] * 32'h029) >> 8) + ((mcu[6][2] * 32'h01b) >> 8) + ((mcu[6][3] * 32'h009) >> 8) + ((mcu[6][4] * -32'h009) >> 8) + ((mcu[6][5] * -32'h01b) >> 8) + ((mcu[6][6] * -32'h029) >> 8) + ((mcu[6][7] * -32'h030) >> 8) + ((mcu[7][0] * -32'h0d0) >> 8) + ((mcu[7][1] * -32'h0b0) >> 8) + ((mcu[7][2] * -32'h076) >> 8) + ((mcu[7][3] * -32'h029) >> 8) + ((mcu[7][4] * 32'h029) >> 8) + ((mcu[7][5] * 32'h076) >> 8) + ((mcu[7][6] * 32'h0b0) >> 8) + ((mcu[7][7] * 32'h0d0) >> 8);
	wire[63:0] cos32_term = ((mcu[0][0] * 32'h0c4) >> 8) + ((mcu[0][1] * 32'h051) >> 8) + ((mcu[0][2] * -32'h051) >> 8) + ((mcu[0][3] * -32'h0c4) >> 8) + ((mcu[0][4] * -32'h0c4) >> 8) + ((mcu[0][5] * -32'h051) >> 8) + ((mcu[0][6] * 32'h051) >> 8) + ((mcu[0][7] * 32'h0c4) >> 8) + ((mcu[1][0] * -32'h02e) >> 8) + ((mcu[1][1] * -32'h013) >> 8) + ((mcu[1][2] * 32'h013) >> 8) + ((mcu[1][3] * 32'h02e) >> 8) + ((mcu[1][4] * 32'h02e) >> 8) + ((mcu[1][5] * 32'h013) >> 8) + ((mcu[1][6] * -32'h013) >> 8) + ((mcu[1][7] * -32'h02e) >> 8) + ((mcu[2][0] * -32'h0e7) >> 8) + ((mcu[2][1] * -32'h060) >> 8) + ((mcu[2][2] * 32'h060) >> 8) + ((mcu[2][3] * 32'h0e7) >> 8) + ((mcu[2][4] * 32'h0e7) >> 8) + ((mcu[2][5] * 32'h060) >> 8) + ((mcu[2][6] * -32'h060) >> 8) + ((mcu[2][7] * -32'h0e7) >> 8) + ((mcu[3][0] * -32'h083) >> 8) + ((mcu[3][1] * -32'h036) >> 8) + ((mcu[3][2] * 32'h036) >> 8) + ((mcu[3][3] * 32'h083) >> 8) + ((mcu[3][4] * 32'h083) >> 8) + ((mcu[3][5] * 32'h036) >> 8) + ((mcu[3][6] * -32'h036) >> 8) + ((mcu[3][7] * -32'h083) >> 8) + ((mcu[4][0] * 32'h083) >> 8) + ((mcu[4][1] * 32'h036) >> 8) + ((mcu[4][2] * -32'h036) >> 8) + ((mcu[4][3] * -32'h083) >> 8) + ((mcu[4][4] * -32'h083) >> 8) + ((mcu[4][5] * -32'h036) >> 8) + ((mcu[4][6] * 32'h036) >> 8) + ((mcu[4][7] * 32'h083) >> 8) + ((mcu[5][0] * 32'h0e7) >> 8) + ((mcu[5][1] * 32'h060) >> 8) + ((mcu[5][2] * -32'h060) >> 8) + ((mcu[5][3] * -32'h0e7) >> 8) + ((mcu[5][4] * -32'h0e7) >> 8) + ((mcu[5][5] * -32'h060) >> 8) + ((mcu[5][6] * 32'h060) >> 8) + ((mcu[5][7] * 32'h0e7) >> 8) + ((mcu[6][0] * 32'h02e) >> 8) + ((mcu[6][1] * 32'h013) >> 8) + ((mcu[6][2] * -32'h013) >> 8) + ((mcu[6][3] * -32'h02e) >> 8) + ((mcu[6][4] * -32'h02e) >> 8) + ((mcu[6][5] * -32'h013) >> 8) + ((mcu[6][6] * 32'h013) >> 8) + ((mcu[6][7] * 32'h02e) >> 8) + ((mcu[7][0] * -32'h0c4) >> 8) + ((mcu[7][1] * -32'h051) >> 8) + ((mcu[7][2] * 32'h051) >> 8) + ((mcu[7][3] * 32'h0c4) >> 8) + ((mcu[7][4] * 32'h0c4) >> 8) + ((mcu[7][5] * 32'h051) >> 8) + ((mcu[7][6] * -32'h051) >> 8) + ((mcu[7][7] * -32'h0c4) >> 8);
	wire[63:0] cos33_term = ((mcu[0][0] * 32'h0b0) >> 8) + ((mcu[0][1] * -32'h029) >> 8) + ((mcu[0][2] * -32'h0d0) >> 8) + ((mcu[0][3] * -32'h076) >> 8) + ((mcu[0][4] * 32'h076) >> 8) + ((mcu[0][5] * 32'h0d0) >> 8) + ((mcu[0][6] * 32'h029) >> 8) + ((mcu[0][7] * -32'h0b0) >> 8) + ((mcu[1][0] * -32'h029) >> 8) + ((mcu[1][1] * 32'h009) >> 8) + ((mcu[1][2] * 32'h030) >> 8) + ((mcu[1][3] * 32'h01b) >> 8) + ((mcu[1][4] * -32'h01b) >> 8) + ((mcu[1][5] * -32'h030) >> 8) + ((mcu[1][6] * -32'h009) >> 8) + ((mcu[1][7] * 32'h029) >> 8) + ((mcu[2][0] * -32'h0d0) >> 8) + ((mcu[2][1] * 32'h030) >> 8) + ((mcu[2][2] * 32'h0f6) >> 8) + ((mcu[2][3] * 32'h08b) >> 8) + ((mcu[2][4] * -32'h08b) >> 8) + ((mcu[2][5] * -32'h0f6) >> 8) + ((mcu[2][6] * -32'h030) >> 8) + ((mcu[2][7] * 32'h0d0) >> 8) + ((mcu[3][0] * -32'h076) >> 8) + ((mcu[3][1] * 32'h01b) >> 8) + ((mcu[3][2] * 32'h08b) >> 8) + ((mcu[3][3] * 32'h04f) >> 8) + ((mcu[3][4] * -32'h04f) >> 8) + ((mcu[3][5] * -32'h08b) >> 8) + ((mcu[3][6] * -32'h01b) >> 8) + ((mcu[3][7] * 32'h076) >> 8) + ((mcu[4][0] * 32'h076) >> 8) + ((mcu[4][1] * -32'h01b) >> 8) + ((mcu[4][2] * -32'h08b) >> 8) + ((mcu[4][3] * -32'h04f) >> 8) + ((mcu[4][4] * 32'h04f) >> 8) + ((mcu[4][5] * 32'h08b) >> 8) + ((mcu[4][6] * 32'h01b) >> 8) + ((mcu[4][7] * -32'h076) >> 8) + ((mcu[5][0] * 32'h0d0) >> 8) + ((mcu[5][1] * -32'h030) >> 8) + ((mcu[5][2] * -32'h0f6) >> 8) + ((mcu[5][3] * -32'h08b) >> 8) + ((mcu[5][4] * 32'h08b) >> 8) + ((mcu[5][5] * 32'h0f6) >> 8) + ((mcu[5][6] * 32'h030) >> 8) + ((mcu[5][7] * -32'h0d0) >> 8) + ((mcu[6][0] * 32'h029) >> 8) + ((mcu[6][1] * -32'h009) >> 8) + ((mcu[6][2] * -32'h030) >> 8) + ((mcu[6][3] * -32'h01b) >> 8) + ((mcu[6][4] * 32'h01b) >> 8) + ((mcu[6][5] * 32'h030) >> 8) + ((mcu[6][6] * 32'h009) >> 8) + ((mcu[6][7] * -32'h029) >> 8) + ((mcu[7][0] * -32'h0b0) >> 8) + ((mcu[7][1] * 32'h029) >> 8) + ((mcu[7][2] * 32'h0d0) >> 8) + ((mcu[7][3] * 32'h076) >> 8) + ((mcu[7][4] * -32'h076) >> 8) + ((mcu[7][5] * -32'h0d0) >> 8) + ((mcu[7][6] * -32'h029) >> 8) + ((mcu[7][7] * 32'h0b0) >> 8);
	wire[63:0] cos34_term = ((mcu[0][0] * 32'h096) >> 8) + ((mcu[0][1] * -32'h096) >> 8) + ((mcu[0][2] * -32'h096) >> 8) + ((mcu[0][3] * 32'h096) >> 8) + ((mcu[0][4] * 32'h096) >> 8) + ((mcu[0][5] * -32'h096) >> 8) + ((mcu[0][6] * -32'h096) >> 8) + ((mcu[0][7] * 32'h096) >> 8) + ((mcu[1][0] * -32'h023) >> 8) + ((mcu[1][1] * 32'h023) >> 8) + ((mcu[1][2] * 32'h023) >> 8) + ((mcu[1][3] * -32'h023) >> 8) + ((mcu[1][4] * -32'h023) >> 8) + ((mcu[1][5] * 32'h023) >> 8) + ((mcu[1][6] * 32'h023) >> 8) + ((mcu[1][7] * -32'h023) >> 8) + ((mcu[2][0] * -32'h0b1) >> 8) + ((mcu[2][1] * 32'h0b1) >> 8) + ((mcu[2][2] * 32'h0b1) >> 8) + ((mcu[2][3] * -32'h0b1) >> 8) + ((mcu[2][4] * -32'h0b1) >> 8) + ((mcu[2][5] * 32'h0b1) >> 8) + ((mcu[2][6] * 32'h0b1) >> 8) + ((mcu[2][7] * -32'h0b1) >> 8) + ((mcu[3][0] * -32'h064) >> 8) + ((mcu[3][1] * 32'h064) >> 8) + ((mcu[3][2] * 32'h064) >> 8) + ((mcu[3][3] * -32'h064) >> 8) + ((mcu[3][4] * -32'h064) >> 8) + ((mcu[3][5] * 32'h064) >> 8) + ((mcu[3][6] * 32'h064) >> 8) + ((mcu[3][7] * -32'h064) >> 8) + ((mcu[4][0] * 32'h064) >> 8) + ((mcu[4][1] * -32'h064) >> 8) + ((mcu[4][2] * -32'h064) >> 8) + ((mcu[4][3] * 32'h064) >> 8) + ((mcu[4][4] * 32'h064) >> 8) + ((mcu[4][5] * -32'h064) >> 8) + ((mcu[4][6] * -32'h064) >> 8) + ((mcu[4][7] * 32'h064) >> 8) + ((mcu[5][0] * 32'h0b1) >> 8) + ((mcu[5][1] * -32'h0b1) >> 8) + ((mcu[5][2] * -32'h0b1) >> 8) + ((mcu[5][3] * 32'h0b1) >> 8) + ((mcu[5][4] * 32'h0b1) >> 8) + ((mcu[5][5] * -32'h0b1) >> 8) + ((mcu[5][6] * -32'h0b1) >> 8) + ((mcu[5][7] * 32'h0b1) >> 8) + ((mcu[6][0] * 32'h023) >> 8) + ((mcu[6][1] * -32'h023) >> 8) + ((mcu[6][2] * -32'h023) >> 8) + ((mcu[6][3] * 32'h023) >> 8) + ((mcu[6][4] * 32'h023) >> 8) + ((mcu[6][5] * -32'h023) >> 8) + ((mcu[6][6] * -32'h023) >> 8) + ((mcu[6][7] * 32'h023) >> 8) + ((mcu[7][0] * -32'h096) >> 8) + ((mcu[7][1] * 32'h096) >> 8) + ((mcu[7][2] * 32'h096) >> 8) + ((mcu[7][3] * -32'h096) >> 8) + ((mcu[7][4] * -32'h096) >> 8) + ((mcu[7][5] * 32'h096) >> 8) + ((mcu[7][6] * 32'h096) >> 8) + ((mcu[7][7] * -32'h096) >> 8);
	wire[63:0] cos35_term = ((mcu[0][0] * 32'h076) >> 8) + ((mcu[0][1] * -32'h0d0) >> 8) + ((mcu[0][2] * 32'h029) >> 8) + ((mcu[0][3] * 32'h0b0) >> 8) + ((mcu[0][4] * -32'h0b0) >> 8) + ((mcu[0][5] * -32'h029) >> 8) + ((mcu[0][6] * 32'h0d0) >> 8) + ((mcu[0][7] * -32'h076) >> 8) + ((mcu[1][0] * -32'h01b) >> 8) + ((mcu[1][1] * 32'h030) >> 8) + ((mcu[1][2] * -32'h009) >> 8) + ((mcu[1][3] * -32'h029) >> 8) + ((mcu[1][4] * 32'h029) >> 8) + ((mcu[1][5] * 32'h009) >> 8) + ((mcu[1][6] * -32'h030) >> 8) + ((mcu[1][7] * 32'h01b) >> 8) + ((mcu[2][0] * -32'h08b) >> 8) + ((mcu[2][1] * 32'h0f6) >> 8) + ((mcu[2][2] * -32'h030) >> 8) + ((mcu[2][3] * -32'h0d0) >> 8) + ((mcu[2][4] * 32'h0d0) >> 8) + ((mcu[2][5] * 32'h030) >> 8) + ((mcu[2][6] * -32'h0f6) >> 8) + ((mcu[2][7] * 32'h08b) >> 8) + ((mcu[3][0] * -32'h04f) >> 8) + ((mcu[3][1] * 32'h08b) >> 8) + ((mcu[3][2] * -32'h01b) >> 8) + ((mcu[3][3] * -32'h076) >> 8) + ((mcu[3][4] * 32'h076) >> 8) + ((mcu[3][5] * 32'h01b) >> 8) + ((mcu[3][6] * -32'h08b) >> 8) + ((mcu[3][7] * 32'h04f) >> 8) + ((mcu[4][0] * 32'h04f) >> 8) + ((mcu[4][1] * -32'h08b) >> 8) + ((mcu[4][2] * 32'h01b) >> 8) + ((mcu[4][3] * 32'h076) >> 8) + ((mcu[4][4] * -32'h076) >> 8) + ((mcu[4][5] * -32'h01b) >> 8) + ((mcu[4][6] * 32'h08b) >> 8) + ((mcu[4][7] * -32'h04f) >> 8) + ((mcu[5][0] * 32'h08b) >> 8) + ((mcu[5][1] * -32'h0f6) >> 8) + ((mcu[5][2] * 32'h030) >> 8) + ((mcu[5][3] * 32'h0d0) >> 8) + ((mcu[5][4] * -32'h0d0) >> 8) + ((mcu[5][5] * -32'h030) >> 8) + ((mcu[5][6] * 32'h0f6) >> 8) + ((mcu[5][7] * -32'h08b) >> 8) + ((mcu[6][0] * 32'h01b) >> 8) + ((mcu[6][1] * -32'h030) >> 8) + ((mcu[6][2] * 32'h009) >> 8) + ((mcu[6][3] * 32'h029) >> 8) + ((mcu[6][4] * -32'h029) >> 8) + ((mcu[6][5] * -32'h009) >> 8) + ((mcu[6][6] * 32'h030) >> 8) + ((mcu[6][7] * -32'h01b) >> 8) + ((mcu[7][0] * -32'h076) >> 8) + ((mcu[7][1] * 32'h0d0) >> 8) + ((mcu[7][2] * -32'h029) >> 8) + ((mcu[7][3] * -32'h0b0) >> 8) + ((mcu[7][4] * 32'h0b0) >> 8) + ((mcu[7][5] * 32'h029) >> 8) + ((mcu[7][6] * -32'h0d0) >> 8) + ((mcu[7][7] * 32'h076) >> 8);
	wire[63:0] cos36_term = ((mcu[0][0] * 32'h051) >> 8) + ((mcu[0][1] * -32'h0c4) >> 8) + ((mcu[0][2] * 32'h0c4) >> 8) + ((mcu[0][3] * -32'h051) >> 8) + ((mcu[0][4] * -32'h051) >> 8) + ((mcu[0][5] * 32'h0c4) >> 8) + ((mcu[0][6] * -32'h0c4) >> 8) + ((mcu[0][7] * 32'h051) >> 8) + ((mcu[1][0] * -32'h013) >> 8) + ((mcu[1][1] * 32'h02e) >> 8) + ((mcu[1][2] * -32'h02e) >> 8) + ((mcu[1][3] * 32'h013) >> 8) + ((mcu[1][4] * 32'h013) >> 8) + ((mcu[1][5] * -32'h02e) >> 8) + ((mcu[1][6] * 32'h02e) >> 8) + ((mcu[1][7] * -32'h013) >> 8) + ((mcu[2][0] * -32'h060) >> 8) + ((mcu[2][1] * 32'h0e7) >> 8) + ((mcu[2][2] * -32'h0e7) >> 8) + ((mcu[2][3] * 32'h060) >> 8) + ((mcu[2][4] * 32'h060) >> 8) + ((mcu[2][5] * -32'h0e7) >> 8) + ((mcu[2][6] * 32'h0e7) >> 8) + ((mcu[2][7] * -32'h060) >> 8) + ((mcu[3][0] * -32'h036) >> 8) + ((mcu[3][1] * 32'h083) >> 8) + ((mcu[3][2] * -32'h083) >> 8) + ((mcu[3][3] * 32'h036) >> 8) + ((mcu[3][4] * 32'h036) >> 8) + ((mcu[3][5] * -32'h083) >> 8) + ((mcu[3][6] * 32'h083) >> 8) + ((mcu[3][7] * -32'h036) >> 8) + ((mcu[4][0] * 32'h036) >> 8) + ((mcu[4][1] * -32'h083) >> 8) + ((mcu[4][2] * 32'h083) >> 8) + ((mcu[4][3] * -32'h036) >> 8) + ((mcu[4][4] * -32'h036) >> 8) + ((mcu[4][5] * 32'h083) >> 8) + ((mcu[4][6] * -32'h083) >> 8) + ((mcu[4][7] * 32'h036) >> 8) + ((mcu[5][0] * 32'h060) >> 8) + ((mcu[5][1] * -32'h0e7) >> 8) + ((mcu[5][2] * 32'h0e7) >> 8) + ((mcu[5][3] * -32'h060) >> 8) + ((mcu[5][4] * -32'h060) >> 8) + ((mcu[5][5] * 32'h0e7) >> 8) + ((mcu[5][6] * -32'h0e7) >> 8) + ((mcu[5][7] * 32'h060) >> 8) + ((mcu[6][0] * 32'h013) >> 8) + ((mcu[6][1] * -32'h02e) >> 8) + ((mcu[6][2] * 32'h02e) >> 8) + ((mcu[6][3] * -32'h013) >> 8) + ((mcu[6][4] * -32'h013) >> 8) + ((mcu[6][5] * 32'h02e) >> 8) + ((mcu[6][6] * -32'h02e) >> 8) + ((mcu[6][7] * 32'h013) >> 8) + ((mcu[7][0] * -32'h051) >> 8) + ((mcu[7][1] * 32'h0c4) >> 8) + ((mcu[7][2] * -32'h0c4) >> 8) + ((mcu[7][3] * 32'h051) >> 8) + ((mcu[7][4] * 32'h051) >> 8) + ((mcu[7][5] * -32'h0c4) >> 8) + ((mcu[7][6] * 32'h0c4) >> 8) + ((mcu[7][7] * -32'h051) >> 8);
	wire[63:0] cos37_term = ((mcu[0][0] * 32'h029) >> 8) + ((mcu[0][1] * -32'h076) >> 8) + ((mcu[0][2] * 32'h0b0) >> 8) + ((mcu[0][3] * -32'h0d0) >> 8) + ((mcu[0][4] * 32'h0d0) >> 8) + ((mcu[0][5] * -32'h0b0) >> 8) + ((mcu[0][6] * 32'h076) >> 8) + ((mcu[0][7] * -32'h029) >> 8) + ((mcu[1][0] * -32'h009) >> 8) + ((mcu[1][1] * 32'h01b) >> 8) + ((mcu[1][2] * -32'h029) >> 8) + ((mcu[1][3] * 32'h030) >> 8) + ((mcu[1][4] * -32'h030) >> 8) + ((mcu[1][5] * 32'h029) >> 8) + ((mcu[1][6] * -32'h01b) >> 8) + ((mcu[1][7] * 32'h009) >> 8) + ((mcu[2][0] * -32'h030) >> 8) + ((mcu[2][1] * 32'h08b) >> 8) + ((mcu[2][2] * -32'h0d0) >> 8) + ((mcu[2][3] * 32'h0f6) >> 8) + ((mcu[2][4] * -32'h0f6) >> 8) + ((mcu[2][5] * 32'h0d0) >> 8) + ((mcu[2][6] * -32'h08b) >> 8) + ((mcu[2][7] * 32'h030) >> 8) + ((mcu[3][0] * -32'h01b) >> 8) + ((mcu[3][1] * 32'h04f) >> 8) + ((mcu[3][2] * -32'h076) >> 8) + ((mcu[3][3] * 32'h08b) >> 8) + ((mcu[3][4] * -32'h08b) >> 8) + ((mcu[3][5] * 32'h076) >> 8) + ((mcu[3][6] * -32'h04f) >> 8) + ((mcu[3][7] * 32'h01b) >> 8) + ((mcu[4][0] * 32'h01b) >> 8) + ((mcu[4][1] * -32'h04f) >> 8) + ((mcu[4][2] * 32'h076) >> 8) + ((mcu[4][3] * -32'h08b) >> 8) + ((mcu[4][4] * 32'h08b) >> 8) + ((mcu[4][5] * -32'h076) >> 8) + ((mcu[4][6] * 32'h04f) >> 8) + ((mcu[4][7] * -32'h01b) >> 8) + ((mcu[5][0] * 32'h030) >> 8) + ((mcu[5][1] * -32'h08b) >> 8) + ((mcu[5][2] * 32'h0d0) >> 8) + ((mcu[5][3] * -32'h0f6) >> 8) + ((mcu[5][4] * 32'h0f6) >> 8) + ((mcu[5][5] * -32'h0d0) >> 8) + ((mcu[5][6] * 32'h08b) >> 8) + ((mcu[5][7] * -32'h030) >> 8) + ((mcu[6][0] * 32'h009) >> 8) + ((mcu[6][1] * -32'h01b) >> 8) + ((mcu[6][2] * 32'h029) >> 8) + ((mcu[6][3] * -32'h030) >> 8) + ((mcu[6][4] * 32'h030) >> 8) + ((mcu[6][5] * -32'h029) >> 8) + ((mcu[6][6] * 32'h01b) >> 8) + ((mcu[6][7] * -32'h009) >> 8) + ((mcu[7][0] * -32'h029) >> 8) + ((mcu[7][1] * 32'h076) >> 8) + ((mcu[7][2] * -32'h0b0) >> 8) + ((mcu[7][3] * 32'h0d0) >> 8) + ((mcu[7][4] * -32'h0d0) >> 8) + ((mcu[7][5] * 32'h0b0) >> 8) + ((mcu[7][6] * -32'h076) >> 8) + ((mcu[7][7] * 32'h029) >> 8);
	wire[63:0] cos40_term = ((mcu[0][0] * 32'h0b4) >> 8) + ((mcu[0][1] * 32'h0b4) >> 8) + ((mcu[0][2] * 32'h0b4) >> 8) + ((mcu[0][3] * 32'h0b4) >> 8) + ((mcu[0][4] * 32'h0b4) >> 8) + ((mcu[0][5] * 32'h0b4) >> 8) + ((mcu[0][6] * 32'h0b4) >> 8) + ((mcu[0][7] * 32'h0b4) >> 8) + ((mcu[1][0] * -32'h0b4) >> 8) + ((mcu[1][1] * -32'h0b4) >> 8) + ((mcu[1][2] * -32'h0b4) >> 8) + ((mcu[1][3] * -32'h0b4) >> 8) + ((mcu[1][4] * -32'h0b4) >> 8) + ((mcu[1][5] * -32'h0b4) >> 8) + ((mcu[1][6] * -32'h0b4) >> 8) + ((mcu[1][7] * -32'h0b4) >> 8) + ((mcu[2][0] * -32'h0b4) >> 8) + ((mcu[2][1] * -32'h0b4) >> 8) + ((mcu[2][2] * -32'h0b4) >> 8) + ((mcu[2][3] * -32'h0b4) >> 8) + ((mcu[2][4] * -32'h0b4) >> 8) + ((mcu[2][5] * -32'h0b4) >> 8) + ((mcu[2][6] * -32'h0b4) >> 8) + ((mcu[2][7] * -32'h0b4) >> 8) + ((mcu[3][0] * 32'h0b4) >> 8) + ((mcu[3][1] * 32'h0b4) >> 8) + ((mcu[3][2] * 32'h0b4) >> 8) + ((mcu[3][3] * 32'h0b4) >> 8) + ((mcu[3][4] * 32'h0b4) >> 8) + ((mcu[3][5] * 32'h0b4) >> 8) + ((mcu[3][6] * 32'h0b4) >> 8) + ((mcu[3][7] * 32'h0b4) >> 8) + ((mcu[4][0] * 32'h0b4) >> 8) + ((mcu[4][1] * 32'h0b4) >> 8) + ((mcu[4][2] * 32'h0b4) >> 8) + ((mcu[4][3] * 32'h0b4) >> 8) + ((mcu[4][4] * 32'h0b4) >> 8) + ((mcu[4][5] * 32'h0b4) >> 8) + ((mcu[4][6] * 32'h0b4) >> 8) + ((mcu[4][7] * 32'h0b4) >> 8) + ((mcu[5][0] * -32'h0b4) >> 8) + ((mcu[5][1] * -32'h0b4) >> 8) + ((mcu[5][2] * -32'h0b4) >> 8) + ((mcu[5][3] * -32'h0b4) >> 8) + ((mcu[5][4] * -32'h0b4) >> 8) + ((mcu[5][5] * -32'h0b4) >> 8) + ((mcu[5][6] * -32'h0b4) >> 8) + ((mcu[5][7] * -32'h0b4) >> 8) + ((mcu[6][0] * -32'h0b4) >> 8) + ((mcu[6][1] * -32'h0b4) >> 8) + ((mcu[6][2] * -32'h0b4) >> 8) + ((mcu[6][3] * -32'h0b4) >> 8) + ((mcu[6][4] * -32'h0b4) >> 8) + ((mcu[6][5] * -32'h0b4) >> 8) + ((mcu[6][6] * -32'h0b4) >> 8) + ((mcu[6][7] * -32'h0b4) >> 8) + ((mcu[7][0] * 32'h0b4) >> 8) + ((mcu[7][1] * 32'h0b4) >> 8) + ((mcu[7][2] * 32'h0b4) >> 8) + ((mcu[7][3] * 32'h0b4) >> 8) + ((mcu[7][4] * 32'h0b4) >> 8) + ((mcu[7][5] * 32'h0b4) >> 8) + ((mcu[7][6] * 32'h0b4) >> 8) + ((mcu[7][7] * 32'h0b4) >> 8);
	wire[63:0] cos41_term = ((mcu[0][0] * 32'h0b1) >> 8) + ((mcu[0][1] * 32'h096) >> 8) + ((mcu[0][2] * 32'h064) >> 8) + ((mcu[0][3] * 32'h023) >> 8) + ((mcu[0][4] * -32'h023) >> 8) + ((mcu[0][5] * -32'h064) >> 8) + ((mcu[0][6] * -32'h096) >> 8) + ((mcu[0][7] * -32'h0b1) >> 8) + ((mcu[1][0] * -32'h0b1) >> 8) + ((mcu[1][1] * -32'h096) >> 8) + ((mcu[1][2] * -32'h064) >> 8) + ((mcu[1][3] * -32'h023) >> 8) + ((mcu[1][4] * 32'h023) >> 8) + ((mcu[1][5] * 32'h064) >> 8) + ((mcu[1][6] * 32'h096) >> 8) + ((mcu[1][7] * 32'h0b1) >> 8) + ((mcu[2][0] * -32'h0b1) >> 8) + ((mcu[2][1] * -32'h096) >> 8) + ((mcu[2][2] * -32'h064) >> 8) + ((mcu[2][3] * -32'h023) >> 8) + ((mcu[2][4] * 32'h023) >> 8) + ((mcu[2][5] * 32'h064) >> 8) + ((mcu[2][6] * 32'h096) >> 8) + ((mcu[2][7] * 32'h0b1) >> 8) + ((mcu[3][0] * 32'h0b1) >> 8) + ((mcu[3][1] * 32'h096) >> 8) + ((mcu[3][2] * 32'h064) >> 8) + ((mcu[3][3] * 32'h023) >> 8) + ((mcu[3][4] * -32'h023) >> 8) + ((mcu[3][5] * -32'h064) >> 8) + ((mcu[3][6] * -32'h096) >> 8) + ((mcu[3][7] * -32'h0b1) >> 8) + ((mcu[4][0] * 32'h0b1) >> 8) + ((mcu[4][1] * 32'h096) >> 8) + ((mcu[4][2] * 32'h064) >> 8) + ((mcu[4][3] * 32'h023) >> 8) + ((mcu[4][4] * -32'h023) >> 8) + ((mcu[4][5] * -32'h064) >> 8) + ((mcu[4][6] * -32'h096) >> 8) + ((mcu[4][7] * -32'h0b1) >> 8) + ((mcu[5][0] * -32'h0b1) >> 8) + ((mcu[5][1] * -32'h096) >> 8) + ((mcu[5][2] * -32'h064) >> 8) + ((mcu[5][3] * -32'h023) >> 8) + ((mcu[5][4] * 32'h023) >> 8) + ((mcu[5][5] * 32'h064) >> 8) + ((mcu[5][6] * 32'h096) >> 8) + ((mcu[5][7] * 32'h0b1) >> 8) + ((mcu[6][0] * -32'h0b1) >> 8) + ((mcu[6][1] * -32'h096) >> 8) + ((mcu[6][2] * -32'h064) >> 8) + ((mcu[6][3] * -32'h023) >> 8) + ((mcu[6][4] * 32'h023) >> 8) + ((mcu[6][5] * 32'h064) >> 8) + ((mcu[6][6] * 32'h096) >> 8) + ((mcu[6][7] * 32'h0b1) >> 8) + ((mcu[7][0] * 32'h0b1) >> 8) + ((mcu[7][1] * 32'h096) >> 8) + ((mcu[7][2] * 32'h064) >> 8) + ((mcu[7][3] * 32'h023) >> 8) + ((mcu[7][4] * -32'h023) >> 8) + ((mcu[7][5] * -32'h064) >> 8) + ((mcu[7][6] * -32'h096) >> 8) + ((mcu[7][7] * -32'h0b1) >> 8);
	wire[63:0] cos42_term = ((mcu[0][0] * 32'h0a7) >> 8) + ((mcu[0][1] * 32'h045) >> 8) + ((mcu[0][2] * -32'h045) >> 8) + ((mcu[0][3] * -32'h0a7) >> 8) + ((mcu[0][4] * -32'h0a7) >> 8) + ((mcu[0][5] * -32'h045) >> 8) + ((mcu[0][6] * 32'h045) >> 8) + ((mcu[0][7] * 32'h0a7) >> 8) + ((mcu[1][0] * -32'h0a7) >> 8) + ((mcu[1][1] * -32'h045) >> 8) + ((mcu[1][2] * 32'h045) >> 8) + ((mcu[1][3] * 32'h0a7) >> 8) + ((mcu[1][4] * 32'h0a7) >> 8) + ((mcu[1][5] * 32'h045) >> 8) + ((mcu[1][6] * -32'h045) >> 8) + ((mcu[1][7] * -32'h0a7) >> 8) + ((mcu[2][0] * -32'h0a7) >> 8) + ((mcu[2][1] * -32'h045) >> 8) + ((mcu[2][2] * 32'h045) >> 8) + ((mcu[2][3] * 32'h0a7) >> 8) + ((mcu[2][4] * 32'h0a7) >> 8) + ((mcu[2][5] * 32'h045) >> 8) + ((mcu[2][6] * -32'h045) >> 8) + ((mcu[2][7] * -32'h0a7) >> 8) + ((mcu[3][0] * 32'h0a7) >> 8) + ((mcu[3][1] * 32'h045) >> 8) + ((mcu[3][2] * -32'h045) >> 8) + ((mcu[3][3] * -32'h0a7) >> 8) + ((mcu[3][4] * -32'h0a7) >> 8) + ((mcu[3][5] * -32'h045) >> 8) + ((mcu[3][6] * 32'h045) >> 8) + ((mcu[3][7] * 32'h0a7) >> 8) + ((mcu[4][0] * 32'h0a7) >> 8) + ((mcu[4][1] * 32'h045) >> 8) + ((mcu[4][2] * -32'h045) >> 8) + ((mcu[4][3] * -32'h0a7) >> 8) + ((mcu[4][4] * -32'h0a7) >> 8) + ((mcu[4][5] * -32'h045) >> 8) + ((mcu[4][6] * 32'h045) >> 8) + ((mcu[4][7] * 32'h0a7) >> 8) + ((mcu[5][0] * -32'h0a7) >> 8) + ((mcu[5][1] * -32'h045) >> 8) + ((mcu[5][2] * 32'h045) >> 8) + ((mcu[5][3] * 32'h0a7) >> 8) + ((mcu[5][4] * 32'h0a7) >> 8) + ((mcu[5][5] * 32'h045) >> 8) + ((mcu[5][6] * -32'h045) >> 8) + ((mcu[5][7] * -32'h0a7) >> 8) + ((mcu[6][0] * -32'h0a7) >> 8) + ((mcu[6][1] * -32'h045) >> 8) + ((mcu[6][2] * 32'h045) >> 8) + ((mcu[6][3] * 32'h0a7) >> 8) + ((mcu[6][4] * 32'h0a7) >> 8) + ((mcu[6][5] * 32'h045) >> 8) + ((mcu[6][6] * -32'h045) >> 8) + ((mcu[6][7] * -32'h0a7) >> 8) + ((mcu[7][0] * 32'h0a7) >> 8) + ((mcu[7][1] * 32'h045) >> 8) + ((mcu[7][2] * -32'h045) >> 8) + ((mcu[7][3] * -32'h0a7) >> 8) + ((mcu[7][4] * -32'h0a7) >> 8) + ((mcu[7][5] * -32'h045) >> 8) + ((mcu[7][6] * 32'h045) >> 8) + ((mcu[7][7] * 32'h0a7) >> 8);
	wire[63:0] cos43_term = ((mcu[0][0] * 32'h096) >> 8) + ((mcu[0][1] * -32'h023) >> 8) + ((mcu[0][2] * -32'h0b1) >> 8) + ((mcu[0][3] * -32'h064) >> 8) + ((mcu[0][4] * 32'h064) >> 8) + ((mcu[0][5] * 32'h0b1) >> 8) + ((mcu[0][6] * 32'h023) >> 8) + ((mcu[0][7] * -32'h096) >> 8) + ((mcu[1][0] * -32'h096) >> 8) + ((mcu[1][1] * 32'h023) >> 8) + ((mcu[1][2] * 32'h0b1) >> 8) + ((mcu[1][3] * 32'h064) >> 8) + ((mcu[1][4] * -32'h064) >> 8) + ((mcu[1][5] * -32'h0b1) >> 8) + ((mcu[1][6] * -32'h023) >> 8) + ((mcu[1][7] * 32'h096) >> 8) + ((mcu[2][0] * -32'h096) >> 8) + ((mcu[2][1] * 32'h023) >> 8) + ((mcu[2][2] * 32'h0b1) >> 8) + ((mcu[2][3] * 32'h064) >> 8) + ((mcu[2][4] * -32'h064) >> 8) + ((mcu[2][5] * -32'h0b1) >> 8) + ((mcu[2][6] * -32'h023) >> 8) + ((mcu[2][7] * 32'h096) >> 8) + ((mcu[3][0] * 32'h096) >> 8) + ((mcu[3][1] * -32'h023) >> 8) + ((mcu[3][2] * -32'h0b1) >> 8) + ((mcu[3][3] * -32'h064) >> 8) + ((mcu[3][4] * 32'h064) >> 8) + ((mcu[3][5] * 32'h0b1) >> 8) + ((mcu[3][6] * 32'h023) >> 8) + ((mcu[3][7] * -32'h096) >> 8) + ((mcu[4][0] * 32'h096) >> 8) + ((mcu[4][1] * -32'h023) >> 8) + ((mcu[4][2] * -32'h0b1) >> 8) + ((mcu[4][3] * -32'h064) >> 8) + ((mcu[4][4] * 32'h064) >> 8) + ((mcu[4][5] * 32'h0b1) >> 8) + ((mcu[4][6] * 32'h023) >> 8) + ((mcu[4][7] * -32'h096) >> 8) + ((mcu[5][0] * -32'h096) >> 8) + ((mcu[5][1] * 32'h023) >> 8) + ((mcu[5][2] * 32'h0b1) >> 8) + ((mcu[5][3] * 32'h064) >> 8) + ((mcu[5][4] * -32'h064) >> 8) + ((mcu[5][5] * -32'h0b1) >> 8) + ((mcu[5][6] * -32'h023) >> 8) + ((mcu[5][7] * 32'h096) >> 8) + ((mcu[6][0] * -32'h096) >> 8) + ((mcu[6][1] * 32'h023) >> 8) + ((mcu[6][2] * 32'h0b1) >> 8) + ((mcu[6][3] * 32'h064) >> 8) + ((mcu[6][4] * -32'h064) >> 8) + ((mcu[6][5] * -32'h0b1) >> 8) + ((mcu[6][6] * -32'h023) >> 8) + ((mcu[6][7] * 32'h096) >> 8) + ((mcu[7][0] * 32'h096) >> 8) + ((mcu[7][1] * -32'h023) >> 8) + ((mcu[7][2] * -32'h0b1) >> 8) + ((mcu[7][3] * -32'h064) >> 8) + ((mcu[7][4] * 32'h064) >> 8) + ((mcu[7][5] * 32'h0b1) >> 8) + ((mcu[7][6] * 32'h023) >> 8) + ((mcu[7][7] * -32'h096) >> 8);
	wire[63:0] cos44_term = ((mcu[0][0] * 32'h080) >> 8) + ((mcu[0][1] * -32'h080) >> 8) + ((mcu[0][2] * -32'h080) >> 8) + ((mcu[0][3] * 32'h080) >> 8) + ((mcu[0][4] * 32'h080) >> 8) + ((mcu[0][5] * -32'h080) >> 8) + ((mcu[0][6] * -32'h080) >> 8) + ((mcu[0][7] * 32'h080) >> 8) + ((mcu[1][0] * -32'h080) >> 8) + ((mcu[1][1] * 32'h080) >> 8) + ((mcu[1][2] * 32'h080) >> 8) + ((mcu[1][3] * -32'h080) >> 8) + ((mcu[1][4] * -32'h080) >> 8) + ((mcu[1][5] * 32'h080) >> 8) + ((mcu[1][6] * 32'h080) >> 8) + ((mcu[1][7] * -32'h080) >> 8) + ((mcu[2][0] * -32'h080) >> 8) + ((mcu[2][1] * 32'h080) >> 8) + ((mcu[2][2] * 32'h080) >> 8) + ((mcu[2][3] * -32'h080) >> 8) + ((mcu[2][4] * -32'h080) >> 8) + ((mcu[2][5] * 32'h080) >> 8) + ((mcu[2][6] * 32'h080) >> 8) + ((mcu[2][7] * -32'h080) >> 8) + ((mcu[3][0] * 32'h080) >> 8) + ((mcu[3][1] * -32'h080) >> 8) + ((mcu[3][2] * -32'h080) >> 8) + ((mcu[3][3] * 32'h080) >> 8) + ((mcu[3][4] * 32'h080) >> 8) + ((mcu[3][5] * -32'h080) >> 8) + ((mcu[3][6] * -32'h080) >> 8) + ((mcu[3][7] * 32'h080) >> 8) + ((mcu[4][0] * 32'h080) >> 8) + ((mcu[4][1] * -32'h080) >> 8) + ((mcu[4][2] * -32'h080) >> 8) + ((mcu[4][3] * 32'h080) >> 8) + ((mcu[4][4] * 32'h080) >> 8) + ((mcu[4][5] * -32'h080) >> 8) + ((mcu[4][6] * -32'h080) >> 8) + ((mcu[4][7] * 32'h080) >> 8) + ((mcu[5][0] * -32'h080) >> 8) + ((mcu[5][1] * 32'h080) >> 8) + ((mcu[5][2] * 32'h080) >> 8) + ((mcu[5][3] * -32'h080) >> 8) + ((mcu[5][4] * -32'h080) >> 8) + ((mcu[5][5] * 32'h080) >> 8) + ((mcu[5][6] * 32'h080) >> 8) + ((mcu[5][7] * -32'h080) >> 8) + ((mcu[6][0] * -32'h080) >> 8) + ((mcu[6][1] * 32'h080) >> 8) + ((mcu[6][2] * 32'h080) >> 8) + ((mcu[6][3] * -32'h080) >> 8) + ((mcu[6][4] * -32'h080) >> 8) + ((mcu[6][5] * 32'h080) >> 8) + ((mcu[6][6] * 32'h080) >> 8) + ((mcu[6][7] * -32'h080) >> 8) + ((mcu[7][0] * 32'h080) >> 8) + ((mcu[7][1] * -32'h080) >> 8) + ((mcu[7][2] * -32'h080) >> 8) + ((mcu[7][3] * 32'h080) >> 8) + ((mcu[7][4] * 32'h080) >> 8) + ((mcu[7][5] * -32'h080) >> 8) + ((mcu[7][6] * -32'h080) >> 8) + ((mcu[7][7] * 32'h080) >> 8);
	wire[63:0] cos45_term = ((mcu[0][0] * 32'h064) >> 8) + ((mcu[0][1] * -32'h0b1) >> 8) + ((mcu[0][2] * 32'h023) >> 8) + ((mcu[0][3] * 32'h096) >> 8) + ((mcu[0][4] * -32'h096) >> 8) + ((mcu[0][5] * -32'h023) >> 8) + ((mcu[0][6] * 32'h0b1) >> 8) + ((mcu[0][7] * -32'h064) >> 8) + ((mcu[1][0] * -32'h064) >> 8) + ((mcu[1][1] * 32'h0b1) >> 8) + ((mcu[1][2] * -32'h023) >> 8) + ((mcu[1][3] * -32'h096) >> 8) + ((mcu[1][4] * 32'h096) >> 8) + ((mcu[1][5] * 32'h023) >> 8) + ((mcu[1][6] * -32'h0b1) >> 8) + ((mcu[1][7] * 32'h064) >> 8) + ((mcu[2][0] * -32'h064) >> 8) + ((mcu[2][1] * 32'h0b1) >> 8) + ((mcu[2][2] * -32'h023) >> 8) + ((mcu[2][3] * -32'h096) >> 8) + ((mcu[2][4] * 32'h096) >> 8) + ((mcu[2][5] * 32'h023) >> 8) + ((mcu[2][6] * -32'h0b1) >> 8) + ((mcu[2][7] * 32'h064) >> 8) + ((mcu[3][0] * 32'h064) >> 8) + ((mcu[3][1] * -32'h0b1) >> 8) + ((mcu[3][2] * 32'h023) >> 8) + ((mcu[3][3] * 32'h096) >> 8) + ((mcu[3][4] * -32'h096) >> 8) + ((mcu[3][5] * -32'h023) >> 8) + ((mcu[3][6] * 32'h0b1) >> 8) + ((mcu[3][7] * -32'h064) >> 8) + ((mcu[4][0] * 32'h064) >> 8) + ((mcu[4][1] * -32'h0b1) >> 8) + ((mcu[4][2] * 32'h023) >> 8) + ((mcu[4][3] * 32'h096) >> 8) + ((mcu[4][4] * -32'h096) >> 8) + ((mcu[4][5] * -32'h023) >> 8) + ((mcu[4][6] * 32'h0b1) >> 8) + ((mcu[4][7] * -32'h064) >> 8) + ((mcu[5][0] * -32'h064) >> 8) + ((mcu[5][1] * 32'h0b1) >> 8) + ((mcu[5][2] * -32'h023) >> 8) + ((mcu[5][3] * -32'h096) >> 8) + ((mcu[5][4] * 32'h096) >> 8) + ((mcu[5][5] * 32'h023) >> 8) + ((mcu[5][6] * -32'h0b1) >> 8) + ((mcu[5][7] * 32'h064) >> 8) + ((mcu[6][0] * -32'h064) >> 8) + ((mcu[6][1] * 32'h0b1) >> 8) + ((mcu[6][2] * -32'h023) >> 8) + ((mcu[6][3] * -32'h096) >> 8) + ((mcu[6][4] * 32'h096) >> 8) + ((mcu[6][5] * 32'h023) >> 8) + ((mcu[6][6] * -32'h0b1) >> 8) + ((mcu[6][7] * 32'h064) >> 8) + ((mcu[7][0] * 32'h064) >> 8) + ((mcu[7][1] * -32'h0b1) >> 8) + ((mcu[7][2] * 32'h023) >> 8) + ((mcu[7][3] * 32'h096) >> 8) + ((mcu[7][4] * -32'h096) >> 8) + ((mcu[7][5] * -32'h023) >> 8) + ((mcu[7][6] * 32'h0b1) >> 8) + ((mcu[7][7] * -32'h064) >> 8);
	wire[63:0] cos46_term = ((mcu[0][0] * 32'h045) >> 8) + ((mcu[0][1] * -32'h0a7) >> 8) + ((mcu[0][2] * 32'h0a7) >> 8) + ((mcu[0][3] * -32'h045) >> 8) + ((mcu[0][4] * -32'h045) >> 8) + ((mcu[0][5] * 32'h0a7) >> 8) + ((mcu[0][6] * -32'h0a7) >> 8) + ((mcu[0][7] * 32'h045) >> 8) + ((mcu[1][0] * -32'h045) >> 8) + ((mcu[1][1] * 32'h0a7) >> 8) + ((mcu[1][2] * -32'h0a7) >> 8) + ((mcu[1][3] * 32'h045) >> 8) + ((mcu[1][4] * 32'h045) >> 8) + ((mcu[1][5] * -32'h0a7) >> 8) + ((mcu[1][6] * 32'h0a7) >> 8) + ((mcu[1][7] * -32'h045) >> 8) + ((mcu[2][0] * -32'h045) >> 8) + ((mcu[2][1] * 32'h0a7) >> 8) + ((mcu[2][2] * -32'h0a7) >> 8) + ((mcu[2][3] * 32'h045) >> 8) + ((mcu[2][4] * 32'h045) >> 8) + ((mcu[2][5] * -32'h0a7) >> 8) + ((mcu[2][6] * 32'h0a7) >> 8) + ((mcu[2][7] * -32'h045) >> 8) + ((mcu[3][0] * 32'h045) >> 8) + ((mcu[3][1] * -32'h0a7) >> 8) + ((mcu[3][2] * 32'h0a7) >> 8) + ((mcu[3][3] * -32'h045) >> 8) + ((mcu[3][4] * -32'h045) >> 8) + ((mcu[3][5] * 32'h0a7) >> 8) + ((mcu[3][6] * -32'h0a7) >> 8) + ((mcu[3][7] * 32'h045) >> 8) + ((mcu[4][0] * 32'h045) >> 8) + ((mcu[4][1] * -32'h0a7) >> 8) + ((mcu[4][2] * 32'h0a7) >> 8) + ((mcu[4][3] * -32'h045) >> 8) + ((mcu[4][4] * -32'h045) >> 8) + ((mcu[4][5] * 32'h0a7) >> 8) + ((mcu[4][6] * -32'h0a7) >> 8) + ((mcu[4][7] * 32'h045) >> 8) + ((mcu[5][0] * -32'h045) >> 8) + ((mcu[5][1] * 32'h0a7) >> 8) + ((mcu[5][2] * -32'h0a7) >> 8) + ((mcu[5][3] * 32'h045) >> 8) + ((mcu[5][4] * 32'h045) >> 8) + ((mcu[5][5] * -32'h0a7) >> 8) + ((mcu[5][6] * 32'h0a7) >> 8) + ((mcu[5][7] * -32'h045) >> 8) + ((mcu[6][0] * -32'h045) >> 8) + ((mcu[6][1] * 32'h0a7) >> 8) + ((mcu[6][2] * -32'h0a7) >> 8) + ((mcu[6][3] * 32'h045) >> 8) + ((mcu[6][4] * 32'h045) >> 8) + ((mcu[6][5] * -32'h0a7) >> 8) + ((mcu[6][6] * 32'h0a7) >> 8) + ((mcu[6][7] * -32'h045) >> 8) + ((mcu[7][0] * 32'h045) >> 8) + ((mcu[7][1] * -32'h0a7) >> 8) + ((mcu[7][2] * 32'h0a7) >> 8) + ((mcu[7][3] * -32'h045) >> 8) + ((mcu[7][4] * -32'h045) >> 8) + ((mcu[7][5] * 32'h0a7) >> 8) + ((mcu[7][6] * -32'h0a7) >> 8) + ((mcu[7][7] * 32'h045) >> 8);
	wire[63:0] cos47_term = ((mcu[0][0] * 32'h023) >> 8) + ((mcu[0][1] * -32'h064) >> 8) + ((mcu[0][2] * 32'h096) >> 8) + ((mcu[0][3] * -32'h0b1) >> 8) + ((mcu[0][4] * 32'h0b1) >> 8) + ((mcu[0][5] * -32'h096) >> 8) + ((mcu[0][6] * 32'h064) >> 8) + ((mcu[0][7] * -32'h023) >> 8) + ((mcu[1][0] * -32'h023) >> 8) + ((mcu[1][1] * 32'h064) >> 8) + ((mcu[1][2] * -32'h096) >> 8) + ((mcu[1][3] * 32'h0b1) >> 8) + ((mcu[1][4] * -32'h0b1) >> 8) + ((mcu[1][5] * 32'h096) >> 8) + ((mcu[1][6] * -32'h064) >> 8) + ((mcu[1][7] * 32'h023) >> 8) + ((mcu[2][0] * -32'h023) >> 8) + ((mcu[2][1] * 32'h064) >> 8) + ((mcu[2][2] * -32'h096) >> 8) + ((mcu[2][3] * 32'h0b1) >> 8) + ((mcu[2][4] * -32'h0b1) >> 8) + ((mcu[2][5] * 32'h096) >> 8) + ((mcu[2][6] * -32'h064) >> 8) + ((mcu[2][7] * 32'h023) >> 8) + ((mcu[3][0] * 32'h023) >> 8) + ((mcu[3][1] * -32'h064) >> 8) + ((mcu[3][2] * 32'h096) >> 8) + ((mcu[3][3] * -32'h0b1) >> 8) + ((mcu[3][4] * 32'h0b1) >> 8) + ((mcu[3][5] * -32'h096) >> 8) + ((mcu[3][6] * 32'h064) >> 8) + ((mcu[3][7] * -32'h023) >> 8) + ((mcu[4][0] * 32'h023) >> 8) + ((mcu[4][1] * -32'h064) >> 8) + ((mcu[4][2] * 32'h096) >> 8) + ((mcu[4][3] * -32'h0b1) >> 8) + ((mcu[4][4] * 32'h0b1) >> 8) + ((mcu[4][5] * -32'h096) >> 8) + ((mcu[4][6] * 32'h064) >> 8) + ((mcu[4][7] * -32'h023) >> 8) + ((mcu[5][0] * -32'h023) >> 8) + ((mcu[5][1] * 32'h064) >> 8) + ((mcu[5][2] * -32'h096) >> 8) + ((mcu[5][3] * 32'h0b1) >> 8) + ((mcu[5][4] * -32'h0b1) >> 8) + ((mcu[5][5] * 32'h096) >> 8) + ((mcu[5][6] * -32'h064) >> 8) + ((mcu[5][7] * 32'h023) >> 8) + ((mcu[6][0] * -32'h023) >> 8) + ((mcu[6][1] * 32'h064) >> 8) + ((mcu[6][2] * -32'h096) >> 8) + ((mcu[6][3] * 32'h0b1) >> 8) + ((mcu[6][4] * -32'h0b1) >> 8) + ((mcu[6][5] * 32'h096) >> 8) + ((mcu[6][6] * -32'h064) >> 8) + ((mcu[6][7] * 32'h023) >> 8) + ((mcu[7][0] * 32'h023) >> 8) + ((mcu[7][1] * -32'h064) >> 8) + ((mcu[7][2] * 32'h096) >> 8) + ((mcu[7][3] * -32'h0b1) >> 8) + ((mcu[7][4] * 32'h0b1) >> 8) + ((mcu[7][5] * -32'h096) >> 8) + ((mcu[7][6] * 32'h064) >> 8) + ((mcu[7][7] * -32'h023) >> 8);
	wire[63:0] cos50_term = ((mcu[0][0] * 32'h08e) >> 8) + ((mcu[0][1] * 32'h08e) >> 8) + ((mcu[0][2] * 32'h08e) >> 8) + ((mcu[0][3] * 32'h08e) >> 8) + ((mcu[0][4] * 32'h08e) >> 8) + ((mcu[0][5] * 32'h08e) >> 8) + ((mcu[0][6] * 32'h08e) >> 8) + ((mcu[0][7] * 32'h08e) >> 8) + ((mcu[1][0] * -32'h0fb) >> 8) + ((mcu[1][1] * -32'h0fb) >> 8) + ((mcu[1][2] * -32'h0fb) >> 8) + ((mcu[1][3] * -32'h0fb) >> 8) + ((mcu[1][4] * -32'h0fb) >> 8) + ((mcu[1][5] * -32'h0fb) >> 8) + ((mcu[1][6] * -32'h0fb) >> 8) + ((mcu[1][7] * -32'h0fb) >> 8) + ((mcu[2][0] * 32'h031) >> 8) + ((mcu[2][1] * 32'h031) >> 8) + ((mcu[2][2] * 32'h031) >> 8) + ((mcu[2][3] * 32'h031) >> 8) + ((mcu[2][4] * 32'h031) >> 8) + ((mcu[2][5] * 32'h031) >> 8) + ((mcu[2][6] * 32'h031) >> 8) + ((mcu[2][7] * 32'h031) >> 8) + ((mcu[3][0] * 32'h0d4) >> 8) + ((mcu[3][1] * 32'h0d4) >> 8) + ((mcu[3][2] * 32'h0d4) >> 8) + ((mcu[3][3] * 32'h0d4) >> 8) + ((mcu[3][4] * 32'h0d4) >> 8) + ((mcu[3][5] * 32'h0d4) >> 8) + ((mcu[3][6] * 32'h0d4) >> 8) + ((mcu[3][7] * 32'h0d4) >> 8) + ((mcu[4][0] * -32'h0d4) >> 8) + ((mcu[4][1] * -32'h0d4) >> 8) + ((mcu[4][2] * -32'h0d4) >> 8) + ((mcu[4][3] * -32'h0d4) >> 8) + ((mcu[4][4] * -32'h0d4) >> 8) + ((mcu[4][5] * -32'h0d4) >> 8) + ((mcu[4][6] * -32'h0d4) >> 8) + ((mcu[4][7] * -32'h0d4) >> 8) + ((mcu[5][0] * -32'h031) >> 8) + ((mcu[5][1] * -32'h031) >> 8) + ((mcu[5][2] * -32'h031) >> 8) + ((mcu[5][3] * -32'h031) >> 8) + ((mcu[5][4] * -32'h031) >> 8) + ((mcu[5][5] * -32'h031) >> 8) + ((mcu[5][6] * -32'h031) >> 8) + ((mcu[5][7] * -32'h031) >> 8) + ((mcu[6][0] * 32'h0fb) >> 8) + ((mcu[6][1] * 32'h0fb) >> 8) + ((mcu[6][2] * 32'h0fb) >> 8) + ((mcu[6][3] * 32'h0fb) >> 8) + ((mcu[6][4] * 32'h0fb) >> 8) + ((mcu[6][5] * 32'h0fb) >> 8) + ((mcu[6][6] * 32'h0fb) >> 8) + ((mcu[6][7] * 32'h0fb) >> 8) + ((mcu[7][0] * -32'h08e) >> 8) + ((mcu[7][1] * -32'h08e) >> 8) + ((mcu[7][2] * -32'h08e) >> 8) + ((mcu[7][3] * -32'h08e) >> 8) + ((mcu[7][4] * -32'h08e) >> 8) + ((mcu[7][5] * -32'h08e) >> 8) + ((mcu[7][6] * -32'h08e) >> 8) + ((mcu[7][7] * -32'h08e) >> 8);
	wire[63:0] cos51_term = ((mcu[0][0] * 32'h08b) >> 8) + ((mcu[0][1] * 32'h076) >> 8) + ((mcu[0][2] * 32'h04f) >> 8) + ((mcu[0][3] * 32'h01b) >> 8) + ((mcu[0][4] * -32'h01b) >> 8) + ((mcu[0][5] * -32'h04f) >> 8) + ((mcu[0][6] * -32'h076) >> 8) + ((mcu[0][7] * -32'h08b) >> 8) + ((mcu[1][0] * -32'h0f6) >> 8) + ((mcu[1][1] * -32'h0d0) >> 8) + ((mcu[1][2] * -32'h08b) >> 8) + ((mcu[1][3] * -32'h030) >> 8) + ((mcu[1][4] * 32'h030) >> 8) + ((mcu[1][5] * 32'h08b) >> 8) + ((mcu[1][6] * 32'h0d0) >> 8) + ((mcu[1][7] * 32'h0f6) >> 8) + ((mcu[2][0] * 32'h030) >> 8) + ((mcu[2][1] * 32'h029) >> 8) + ((mcu[2][2] * 32'h01b) >> 8) + ((mcu[2][3] * 32'h009) >> 8) + ((mcu[2][4] * -32'h009) >> 8) + ((mcu[2][5] * -32'h01b) >> 8) + ((mcu[2][6] * -32'h029) >> 8) + ((mcu[2][7] * -32'h030) >> 8) + ((mcu[3][0] * 32'h0d0) >> 8) + ((mcu[3][1] * 32'h0b0) >> 8) + ((mcu[3][2] * 32'h076) >> 8) + ((mcu[3][3] * 32'h029) >> 8) + ((mcu[3][4] * -32'h029) >> 8) + ((mcu[3][5] * -32'h076) >> 8) + ((mcu[3][6] * -32'h0b0) >> 8) + ((mcu[3][7] * -32'h0d0) >> 8) + ((mcu[4][0] * -32'h0d0) >> 8) + ((mcu[4][1] * -32'h0b0) >> 8) + ((mcu[4][2] * -32'h076) >> 8) + ((mcu[4][3] * -32'h029) >> 8) + ((mcu[4][4] * 32'h029) >> 8) + ((mcu[4][5] * 32'h076) >> 8) + ((mcu[4][6] * 32'h0b0) >> 8) + ((mcu[4][7] * 32'h0d0) >> 8) + ((mcu[5][0] * -32'h030) >> 8) + ((mcu[5][1] * -32'h029) >> 8) + ((mcu[5][2] * -32'h01b) >> 8) + ((mcu[5][3] * -32'h009) >> 8) + ((mcu[5][4] * 32'h009) >> 8) + ((mcu[5][5] * 32'h01b) >> 8) + ((mcu[5][6] * 32'h029) >> 8) + ((mcu[5][7] * 32'h030) >> 8) + ((mcu[6][0] * 32'h0f6) >> 8) + ((mcu[6][1] * 32'h0d0) >> 8) + ((mcu[6][2] * 32'h08b) >> 8) + ((mcu[6][3] * 32'h030) >> 8) + ((mcu[6][4] * -32'h030) >> 8) + ((mcu[6][5] * -32'h08b) >> 8) + ((mcu[6][6] * -32'h0d0) >> 8) + ((mcu[6][7] * -32'h0f6) >> 8) + ((mcu[7][0] * -32'h08b) >> 8) + ((mcu[7][1] * -32'h076) >> 8) + ((mcu[7][2] * -32'h04f) >> 8) + ((mcu[7][3] * -32'h01b) >> 8) + ((mcu[7][4] * 32'h01b) >> 8) + ((mcu[7][5] * 32'h04f) >> 8) + ((mcu[7][6] * 32'h076) >> 8) + ((mcu[7][7] * 32'h08b) >> 8);
	wire[63:0] cos52_term = ((mcu[0][0] * 32'h083) >> 8) + ((mcu[0][1] * 32'h036) >> 8) + ((mcu[0][2] * -32'h036) >> 8) + ((mcu[0][3] * -32'h083) >> 8) + ((mcu[0][4] * -32'h083) >> 8) + ((mcu[0][5] * -32'h036) >> 8) + ((mcu[0][6] * 32'h036) >> 8) + ((mcu[0][7] * 32'h083) >> 8) + ((mcu[1][0] * -32'h0e7) >> 8) + ((mcu[1][1] * -32'h060) >> 8) + ((mcu[1][2] * 32'h060) >> 8) + ((mcu[1][3] * 32'h0e7) >> 8) + ((mcu[1][4] * 32'h0e7) >> 8) + ((mcu[1][5] * 32'h060) >> 8) + ((mcu[1][6] * -32'h060) >> 8) + ((mcu[1][7] * -32'h0e7) >> 8) + ((mcu[2][0] * 32'h02e) >> 8) + ((mcu[2][1] * 32'h013) >> 8) + ((mcu[2][2] * -32'h013) >> 8) + ((mcu[2][3] * -32'h02e) >> 8) + ((mcu[2][4] * -32'h02e) >> 8) + ((mcu[2][5] * -32'h013) >> 8) + ((mcu[2][6] * 32'h013) >> 8) + ((mcu[2][7] * 32'h02e) >> 8) + ((mcu[3][0] * 32'h0c4) >> 8) + ((mcu[3][1] * 32'h051) >> 8) + ((mcu[3][2] * -32'h051) >> 8) + ((mcu[3][3] * -32'h0c4) >> 8) + ((mcu[3][4] * -32'h0c4) >> 8) + ((mcu[3][5] * -32'h051) >> 8) + ((mcu[3][6] * 32'h051) >> 8) + ((mcu[3][7] * 32'h0c4) >> 8) + ((mcu[4][0] * -32'h0c4) >> 8) + ((mcu[4][1] * -32'h051) >> 8) + ((mcu[4][2] * 32'h051) >> 8) + ((mcu[4][3] * 32'h0c4) >> 8) + ((mcu[4][4] * 32'h0c4) >> 8) + ((mcu[4][5] * 32'h051) >> 8) + ((mcu[4][6] * -32'h051) >> 8) + ((mcu[4][7] * -32'h0c4) >> 8) + ((mcu[5][0] * -32'h02e) >> 8) + ((mcu[5][1] * -32'h013) >> 8) + ((mcu[5][2] * 32'h013) >> 8) + ((mcu[5][3] * 32'h02e) >> 8) + ((mcu[5][4] * 32'h02e) >> 8) + ((mcu[5][5] * 32'h013) >> 8) + ((mcu[5][6] * -32'h013) >> 8) + ((mcu[5][7] * -32'h02e) >> 8) + ((mcu[6][0] * 32'h0e7) >> 8) + ((mcu[6][1] * 32'h060) >> 8) + ((mcu[6][2] * -32'h060) >> 8) + ((mcu[6][3] * -32'h0e7) >> 8) + ((mcu[6][4] * -32'h0e7) >> 8) + ((mcu[6][5] * -32'h060) >> 8) + ((mcu[6][6] * 32'h060) >> 8) + ((mcu[6][7] * 32'h0e7) >> 8) + ((mcu[7][0] * -32'h083) >> 8) + ((mcu[7][1] * -32'h036) >> 8) + ((mcu[7][2] * 32'h036) >> 8) + ((mcu[7][3] * 32'h083) >> 8) + ((mcu[7][4] * 32'h083) >> 8) + ((mcu[7][5] * 32'h036) >> 8) + ((mcu[7][6] * -32'h036) >> 8) + ((mcu[7][7] * -32'h083) >> 8);
	wire[63:0] cos53_term = ((mcu[0][0] * 32'h076) >> 8) + ((mcu[0][1] * -32'h01b) >> 8) + ((mcu[0][2] * -32'h08b) >> 8) + ((mcu[0][3] * -32'h04f) >> 8) + ((mcu[0][4] * 32'h04f) >> 8) + ((mcu[0][5] * 32'h08b) >> 8) + ((mcu[0][6] * 32'h01b) >> 8) + ((mcu[0][7] * -32'h076) >> 8) + ((mcu[1][0] * -32'h0d0) >> 8) + ((mcu[1][1] * 32'h030) >> 8) + ((mcu[1][2] * 32'h0f6) >> 8) + ((mcu[1][3] * 32'h08b) >> 8) + ((mcu[1][4] * -32'h08b) >> 8) + ((mcu[1][5] * -32'h0f6) >> 8) + ((mcu[1][6] * -32'h030) >> 8) + ((mcu[1][7] * 32'h0d0) >> 8) + ((mcu[2][0] * 32'h029) >> 8) + ((mcu[2][1] * -32'h009) >> 8) + ((mcu[2][2] * -32'h030) >> 8) + ((mcu[2][3] * -32'h01b) >> 8) + ((mcu[2][4] * 32'h01b) >> 8) + ((mcu[2][5] * 32'h030) >> 8) + ((mcu[2][6] * 32'h009) >> 8) + ((mcu[2][7] * -32'h029) >> 8) + ((mcu[3][0] * 32'h0b0) >> 8) + ((mcu[3][1] * -32'h029) >> 8) + ((mcu[3][2] * -32'h0d0) >> 8) + ((mcu[3][3] * -32'h076) >> 8) + ((mcu[3][4] * 32'h076) >> 8) + ((mcu[3][5] * 32'h0d0) >> 8) + ((mcu[3][6] * 32'h029) >> 8) + ((mcu[3][7] * -32'h0b0) >> 8) + ((mcu[4][0] * -32'h0b0) >> 8) + ((mcu[4][1] * 32'h029) >> 8) + ((mcu[4][2] * 32'h0d0) >> 8) + ((mcu[4][3] * 32'h076) >> 8) + ((mcu[4][4] * -32'h076) >> 8) + ((mcu[4][5] * -32'h0d0) >> 8) + ((mcu[4][6] * -32'h029) >> 8) + ((mcu[4][7] * 32'h0b0) >> 8) + ((mcu[5][0] * -32'h029) >> 8) + ((mcu[5][1] * 32'h009) >> 8) + ((mcu[5][2] * 32'h030) >> 8) + ((mcu[5][3] * 32'h01b) >> 8) + ((mcu[5][4] * -32'h01b) >> 8) + ((mcu[5][5] * -32'h030) >> 8) + ((mcu[5][6] * -32'h009) >> 8) + ((mcu[5][7] * 32'h029) >> 8) + ((mcu[6][0] * 32'h0d0) >> 8) + ((mcu[6][1] * -32'h030) >> 8) + ((mcu[6][2] * -32'h0f6) >> 8) + ((mcu[6][3] * -32'h08b) >> 8) + ((mcu[6][4] * 32'h08b) >> 8) + ((mcu[6][5] * 32'h0f6) >> 8) + ((mcu[6][6] * 32'h030) >> 8) + ((mcu[6][7] * -32'h0d0) >> 8) + ((mcu[7][0] * -32'h076) >> 8) + ((mcu[7][1] * 32'h01b) >> 8) + ((mcu[7][2] * 32'h08b) >> 8) + ((mcu[7][3] * 32'h04f) >> 8) + ((mcu[7][4] * -32'h04f) >> 8) + ((mcu[7][5] * -32'h08b) >> 8) + ((mcu[7][6] * -32'h01b) >> 8) + ((mcu[7][7] * 32'h076) >> 8);
	wire[63:0] cos54_term = ((mcu[0][0] * 32'h064) >> 8) + ((mcu[0][1] * -32'h064) >> 8) + ((mcu[0][2] * -32'h064) >> 8) + ((mcu[0][3] * 32'h064) >> 8) + ((mcu[0][4] * 32'h064) >> 8) + ((mcu[0][5] * -32'h064) >> 8) + ((mcu[0][6] * -32'h064) >> 8) + ((mcu[0][7] * 32'h064) >> 8) + ((mcu[1][0] * -32'h0b1) >> 8) + ((mcu[1][1] * 32'h0b1) >> 8) + ((mcu[1][2] * 32'h0b1) >> 8) + ((mcu[1][3] * -32'h0b1) >> 8) + ((mcu[1][4] * -32'h0b1) >> 8) + ((mcu[1][5] * 32'h0b1) >> 8) + ((mcu[1][6] * 32'h0b1) >> 8) + ((mcu[1][7] * -32'h0b1) >> 8) + ((mcu[2][0] * 32'h023) >> 8) + ((mcu[2][1] * -32'h023) >> 8) + ((mcu[2][2] * -32'h023) >> 8) + ((mcu[2][3] * 32'h023) >> 8) + ((mcu[2][4] * 32'h023) >> 8) + ((mcu[2][5] * -32'h023) >> 8) + ((mcu[2][6] * -32'h023) >> 8) + ((mcu[2][7] * 32'h023) >> 8) + ((mcu[3][0] * 32'h096) >> 8) + ((mcu[3][1] * -32'h096) >> 8) + ((mcu[3][2] * -32'h096) >> 8) + ((mcu[3][3] * 32'h096) >> 8) + ((mcu[3][4] * 32'h096) >> 8) + ((mcu[3][5] * -32'h096) >> 8) + ((mcu[3][6] * -32'h096) >> 8) + ((mcu[3][7] * 32'h096) >> 8) + ((mcu[4][0] * -32'h096) >> 8) + ((mcu[4][1] * 32'h096) >> 8) + ((mcu[4][2] * 32'h096) >> 8) + ((mcu[4][3] * -32'h096) >> 8) + ((mcu[4][4] * -32'h096) >> 8) + ((mcu[4][5] * 32'h096) >> 8) + ((mcu[4][6] * 32'h096) >> 8) + ((mcu[4][7] * -32'h096) >> 8) + ((mcu[5][0] * -32'h023) >> 8) + ((mcu[5][1] * 32'h023) >> 8) + ((mcu[5][2] * 32'h023) >> 8) + ((mcu[5][3] * -32'h023) >> 8) + ((mcu[5][4] * -32'h023) >> 8) + ((mcu[5][5] * 32'h023) >> 8) + ((mcu[5][6] * 32'h023) >> 8) + ((mcu[5][7] * -32'h023) >> 8) + ((mcu[6][0] * 32'h0b1) >> 8) + ((mcu[6][1] * -32'h0b1) >> 8) + ((mcu[6][2] * -32'h0b1) >> 8) + ((mcu[6][3] * 32'h0b1) >> 8) + ((mcu[6][4] * 32'h0b1) >> 8) + ((mcu[6][5] * -32'h0b1) >> 8) + ((mcu[6][6] * -32'h0b1) >> 8) + ((mcu[6][7] * 32'h0b1) >> 8) + ((mcu[7][0] * -32'h064) >> 8) + ((mcu[7][1] * 32'h064) >> 8) + ((mcu[7][2] * 32'h064) >> 8) + ((mcu[7][3] * -32'h064) >> 8) + ((mcu[7][4] * -32'h064) >> 8) + ((mcu[7][5] * 32'h064) >> 8) + ((mcu[7][6] * 32'h064) >> 8) + ((mcu[7][7] * -32'h064) >> 8);
	wire[63:0] cos55_term = ((mcu[0][0] * 32'h04f) >> 8) + ((mcu[0][1] * -32'h08b) >> 8) + ((mcu[0][2] * 32'h01b) >> 8) + ((mcu[0][3] * 32'h076) >> 8) + ((mcu[0][4] * -32'h076) >> 8) + ((mcu[0][5] * -32'h01b) >> 8) + ((mcu[0][6] * 32'h08b) >> 8) + ((mcu[0][7] * -32'h04f) >> 8) + ((mcu[1][0] * -32'h08b) >> 8) + ((mcu[1][1] * 32'h0f6) >> 8) + ((mcu[1][2] * -32'h030) >> 8) + ((mcu[1][3] * -32'h0d0) >> 8) + ((mcu[1][4] * 32'h0d0) >> 8) + ((mcu[1][5] * 32'h030) >> 8) + ((mcu[1][6] * -32'h0f6) >> 8) + ((mcu[1][7] * 32'h08b) >> 8) + ((mcu[2][0] * 32'h01b) >> 8) + ((mcu[2][1] * -32'h030) >> 8) + ((mcu[2][2] * 32'h009) >> 8) + ((mcu[2][3] * 32'h029) >> 8) + ((mcu[2][4] * -32'h029) >> 8) + ((mcu[2][5] * -32'h009) >> 8) + ((mcu[2][6] * 32'h030) >> 8) + ((mcu[2][7] * -32'h01b) >> 8) + ((mcu[3][0] * 32'h076) >> 8) + ((mcu[3][1] * -32'h0d0) >> 8) + ((mcu[3][2] * 32'h029) >> 8) + ((mcu[3][3] * 32'h0b0) >> 8) + ((mcu[3][4] * -32'h0b0) >> 8) + ((mcu[3][5] * -32'h029) >> 8) + ((mcu[3][6] * 32'h0d0) >> 8) + ((mcu[3][7] * -32'h076) >> 8) + ((mcu[4][0] * -32'h076) >> 8) + ((mcu[4][1] * 32'h0d0) >> 8) + ((mcu[4][2] * -32'h029) >> 8) + ((mcu[4][3] * -32'h0b0) >> 8) + ((mcu[4][4] * 32'h0b0) >> 8) + ((mcu[4][5] * 32'h029) >> 8) + ((mcu[4][6] * -32'h0d0) >> 8) + ((mcu[4][7] * 32'h076) >> 8) + ((mcu[5][0] * -32'h01b) >> 8) + ((mcu[5][1] * 32'h030) >> 8) + ((mcu[5][2] * -32'h009) >> 8) + ((mcu[5][3] * -32'h029) >> 8) + ((mcu[5][4] * 32'h029) >> 8) + ((mcu[5][5] * 32'h009) >> 8) + ((mcu[5][6] * -32'h030) >> 8) + ((mcu[5][7] * 32'h01b) >> 8) + ((mcu[6][0] * 32'h08b) >> 8) + ((mcu[6][1] * -32'h0f6) >> 8) + ((mcu[6][2] * 32'h030) >> 8) + ((mcu[6][3] * 32'h0d0) >> 8) + ((mcu[6][4] * -32'h0d0) >> 8) + ((mcu[6][5] * -32'h030) >> 8) + ((mcu[6][6] * 32'h0f6) >> 8) + ((mcu[6][7] * -32'h08b) >> 8) + ((mcu[7][0] * -32'h04f) >> 8) + ((mcu[7][1] * 32'h08b) >> 8) + ((mcu[7][2] * -32'h01b) >> 8) + ((mcu[7][3] * -32'h076) >> 8) + ((mcu[7][4] * 32'h076) >> 8) + ((mcu[7][5] * 32'h01b) >> 8) + ((mcu[7][6] * -32'h08b) >> 8) + ((mcu[7][7] * 32'h04f) >> 8);
	wire[63:0] cos56_term = ((mcu[0][0] * 32'h036) >> 8) + ((mcu[0][1] * -32'h083) >> 8) + ((mcu[0][2] * 32'h083) >> 8) + ((mcu[0][3] * -32'h036) >> 8) + ((mcu[0][4] * -32'h036) >> 8) + ((mcu[0][5] * 32'h083) >> 8) + ((mcu[0][6] * -32'h083) >> 8) + ((mcu[0][7] * 32'h036) >> 8) + ((mcu[1][0] * -32'h060) >> 8) + ((mcu[1][1] * 32'h0e7) >> 8) + ((mcu[1][2] * -32'h0e7) >> 8) + ((mcu[1][3] * 32'h060) >> 8) + ((mcu[1][4] * 32'h060) >> 8) + ((mcu[1][5] * -32'h0e7) >> 8) + ((mcu[1][6] * 32'h0e7) >> 8) + ((mcu[1][7] * -32'h060) >> 8) + ((mcu[2][0] * 32'h013) >> 8) + ((mcu[2][1] * -32'h02e) >> 8) + ((mcu[2][2] * 32'h02e) >> 8) + ((mcu[2][3] * -32'h013) >> 8) + ((mcu[2][4] * -32'h013) >> 8) + ((mcu[2][5] * 32'h02e) >> 8) + ((mcu[2][6] * -32'h02e) >> 8) + ((mcu[2][7] * 32'h013) >> 8) + ((mcu[3][0] * 32'h051) >> 8) + ((mcu[3][1] * -32'h0c4) >> 8) + ((mcu[3][2] * 32'h0c4) >> 8) + ((mcu[3][3] * -32'h051) >> 8) + ((mcu[3][4] * -32'h051) >> 8) + ((mcu[3][5] * 32'h0c4) >> 8) + ((mcu[3][6] * -32'h0c4) >> 8) + ((mcu[3][7] * 32'h051) >> 8) + ((mcu[4][0] * -32'h051) >> 8) + ((mcu[4][1] * 32'h0c4) >> 8) + ((mcu[4][2] * -32'h0c4) >> 8) + ((mcu[4][3] * 32'h051) >> 8) + ((mcu[4][4] * 32'h051) >> 8) + ((mcu[4][5] * -32'h0c4) >> 8) + ((mcu[4][6] * 32'h0c4) >> 8) + ((mcu[4][7] * -32'h051) >> 8) + ((mcu[5][0] * -32'h013) >> 8) + ((mcu[5][1] * 32'h02e) >> 8) + ((mcu[5][2] * -32'h02e) >> 8) + ((mcu[5][3] * 32'h013) >> 8) + ((mcu[5][4] * 32'h013) >> 8) + ((mcu[5][5] * -32'h02e) >> 8) + ((mcu[5][6] * 32'h02e) >> 8) + ((mcu[5][7] * -32'h013) >> 8) + ((mcu[6][0] * 32'h060) >> 8) + ((mcu[6][1] * -32'h0e7) >> 8) + ((mcu[6][2] * 32'h0e7) >> 8) + ((mcu[6][3] * -32'h060) >> 8) + ((mcu[6][4] * -32'h060) >> 8) + ((mcu[6][5] * 32'h0e7) >> 8) + ((mcu[6][6] * -32'h0e7) >> 8) + ((mcu[6][7] * 32'h060) >> 8) + ((mcu[7][0] * -32'h036) >> 8) + ((mcu[7][1] * 32'h083) >> 8) + ((mcu[7][2] * -32'h083) >> 8) + ((mcu[7][3] * 32'h036) >> 8) + ((mcu[7][4] * 32'h036) >> 8) + ((mcu[7][5] * -32'h083) >> 8) + ((mcu[7][6] * 32'h083) >> 8) + ((mcu[7][7] * -32'h036) >> 8);
	wire[63:0] cos57_term = ((mcu[0][0] * 32'h01b) >> 8) + ((mcu[0][1] * -32'h04f) >> 8) + ((mcu[0][2] * 32'h076) >> 8) + ((mcu[0][3] * -32'h08b) >> 8) + ((mcu[0][4] * 32'h08b) >> 8) + ((mcu[0][5] * -32'h076) >> 8) + ((mcu[0][6] * 32'h04f) >> 8) + ((mcu[0][7] * -32'h01b) >> 8) + ((mcu[1][0] * -32'h030) >> 8) + ((mcu[1][1] * 32'h08b) >> 8) + ((mcu[1][2] * -32'h0d0) >> 8) + ((mcu[1][3] * 32'h0f6) >> 8) + ((mcu[1][4] * -32'h0f6) >> 8) + ((mcu[1][5] * 32'h0d0) >> 8) + ((mcu[1][6] * -32'h08b) >> 8) + ((mcu[1][7] * 32'h030) >> 8) + ((mcu[2][0] * 32'h009) >> 8) + ((mcu[2][1] * -32'h01b) >> 8) + ((mcu[2][2] * 32'h029) >> 8) + ((mcu[2][3] * -32'h030) >> 8) + ((mcu[2][4] * 32'h030) >> 8) + ((mcu[2][5] * -32'h029) >> 8) + ((mcu[2][6] * 32'h01b) >> 8) + ((mcu[2][7] * -32'h009) >> 8) + ((mcu[3][0] * 32'h029) >> 8) + ((mcu[3][1] * -32'h076) >> 8) + ((mcu[3][2] * 32'h0b0) >> 8) + ((mcu[3][3] * -32'h0d0) >> 8) + ((mcu[3][4] * 32'h0d0) >> 8) + ((mcu[3][5] * -32'h0b0) >> 8) + ((mcu[3][6] * 32'h076) >> 8) + ((mcu[3][7] * -32'h029) >> 8) + ((mcu[4][0] * -32'h029) >> 8) + ((mcu[4][1] * 32'h076) >> 8) + ((mcu[4][2] * -32'h0b0) >> 8) + ((mcu[4][3] * 32'h0d0) >> 8) + ((mcu[4][4] * -32'h0d0) >> 8) + ((mcu[4][5] * 32'h0b0) >> 8) + ((mcu[4][6] * -32'h076) >> 8) + ((mcu[4][7] * 32'h029) >> 8) + ((mcu[5][0] * -32'h009) >> 8) + ((mcu[5][1] * 32'h01b) >> 8) + ((mcu[5][2] * -32'h029) >> 8) + ((mcu[5][3] * 32'h030) >> 8) + ((mcu[5][4] * -32'h030) >> 8) + ((mcu[5][5] * 32'h029) >> 8) + ((mcu[5][6] * -32'h01b) >> 8) + ((mcu[5][7] * 32'h009) >> 8) + ((mcu[6][0] * 32'h030) >> 8) + ((mcu[6][1] * -32'h08b) >> 8) + ((mcu[6][2] * 32'h0d0) >> 8) + ((mcu[6][3] * -32'h0f6) >> 8) + ((mcu[6][4] * 32'h0f6) >> 8) + ((mcu[6][5] * -32'h0d0) >> 8) + ((mcu[6][6] * 32'h08b) >> 8) + ((mcu[6][7] * -32'h030) >> 8) + ((mcu[7][0] * -32'h01b) >> 8) + ((mcu[7][1] * 32'h04f) >> 8) + ((mcu[7][2] * -32'h076) >> 8) + ((mcu[7][3] * 32'h08b) >> 8) + ((mcu[7][4] * -32'h08b) >> 8) + ((mcu[7][5] * 32'h076) >> 8) + ((mcu[7][6] * -32'h04f) >> 8) + ((mcu[7][7] * 32'h01b) >> 8);
	wire[63:0] cos60_term = ((mcu[0][0] * 32'h062) >> 8) + ((mcu[0][1] * 32'h062) >> 8) + ((mcu[0][2] * 32'h062) >> 8) + ((mcu[0][3] * 32'h062) >> 8) + ((mcu[0][4] * 32'h062) >> 8) + ((mcu[0][5] * 32'h062) >> 8) + ((mcu[0][6] * 32'h062) >> 8) + ((mcu[0][7] * 32'h062) >> 8) + ((mcu[1][0] * -32'h0ec) >> 8) + ((mcu[1][1] * -32'h0ec) >> 8) + ((mcu[1][2] * -32'h0ec) >> 8) + ((mcu[1][3] * -32'h0ec) >> 8) + ((mcu[1][4] * -32'h0ec) >> 8) + ((mcu[1][5] * -32'h0ec) >> 8) + ((mcu[1][6] * -32'h0ec) >> 8) + ((mcu[1][7] * -32'h0ec) >> 8) + ((mcu[2][0] * 32'h0ec) >> 8) + ((mcu[2][1] * 32'h0ec) >> 8) + ((mcu[2][2] * 32'h0ec) >> 8) + ((mcu[2][3] * 32'h0ec) >> 8) + ((mcu[2][4] * 32'h0ec) >> 8) + ((mcu[2][5] * 32'h0ec) >> 8) + ((mcu[2][6] * 32'h0ec) >> 8) + ((mcu[2][7] * 32'h0ec) >> 8) + ((mcu[3][0] * -32'h062) >> 8) + ((mcu[3][1] * -32'h062) >> 8) + ((mcu[3][2] * -32'h062) >> 8) + ((mcu[3][3] * -32'h062) >> 8) + ((mcu[3][4] * -32'h062) >> 8) + ((mcu[3][5] * -32'h062) >> 8) + ((mcu[3][6] * -32'h062) >> 8) + ((mcu[3][7] * -32'h062) >> 8) + ((mcu[4][0] * -32'h062) >> 8) + ((mcu[4][1] * -32'h062) >> 8) + ((mcu[4][2] * -32'h062) >> 8) + ((mcu[4][3] * -32'h062) >> 8) + ((mcu[4][4] * -32'h062) >> 8) + ((mcu[4][5] * -32'h062) >> 8) + ((mcu[4][6] * -32'h062) >> 8) + ((mcu[4][7] * -32'h062) >> 8) + ((mcu[5][0] * 32'h0ec) >> 8) + ((mcu[5][1] * 32'h0ec) >> 8) + ((mcu[5][2] * 32'h0ec) >> 8) + ((mcu[5][3] * 32'h0ec) >> 8) + ((mcu[5][4] * 32'h0ec) >> 8) + ((mcu[5][5] * 32'h0ec) >> 8) + ((mcu[5][6] * 32'h0ec) >> 8) + ((mcu[5][7] * 32'h0ec) >> 8) + ((mcu[6][0] * -32'h0ec) >> 8) + ((mcu[6][1] * -32'h0ec) >> 8) + ((mcu[6][2] * -32'h0ec) >> 8) + ((mcu[6][3] * -32'h0ec) >> 8) + ((mcu[6][4] * -32'h0ec) >> 8) + ((mcu[6][5] * -32'h0ec) >> 8) + ((mcu[6][6] * -32'h0ec) >> 8) + ((mcu[6][7] * -32'h0ec) >> 8) + ((mcu[7][0] * 32'h062) >> 8) + ((mcu[7][1] * 32'h062) >> 8) + ((mcu[7][2] * 32'h062) >> 8) + ((mcu[7][3] * 32'h062) >> 8) + ((mcu[7][4] * 32'h062) >> 8) + ((mcu[7][5] * 32'h062) >> 8) + ((mcu[7][6] * 32'h062) >> 8) + ((mcu[7][7] * 32'h062) >> 8);
	wire[63:0] cos61_term = ((mcu[0][0] * 32'h060) >> 8) + ((mcu[0][1] * 32'h051) >> 8) + ((mcu[0][2] * 32'h036) >> 8) + ((mcu[0][3] * 32'h013) >> 8) + ((mcu[0][4] * -32'h013) >> 8) + ((mcu[0][5] * -32'h036) >> 8) + ((mcu[0][6] * -32'h051) >> 8) + ((mcu[0][7] * -32'h060) >> 8) + ((mcu[1][0] * -32'h0e7) >> 8) + ((mcu[1][1] * -32'h0c4) >> 8) + ((mcu[1][2] * -32'h083) >> 8) + ((mcu[1][3] * -32'h02e) >> 8) + ((mcu[1][4] * 32'h02e) >> 8) + ((mcu[1][5] * 32'h083) >> 8) + ((mcu[1][6] * 32'h0c4) >> 8) + ((mcu[1][7] * 32'h0e7) >> 8) + ((mcu[2][0] * 32'h0e7) >> 8) + ((mcu[2][1] * 32'h0c4) >> 8) + ((mcu[2][2] * 32'h083) >> 8) + ((mcu[2][3] * 32'h02e) >> 8) + ((mcu[2][4] * -32'h02e) >> 8) + ((mcu[2][5] * -32'h083) >> 8) + ((mcu[2][6] * -32'h0c4) >> 8) + ((mcu[2][7] * -32'h0e7) >> 8) + ((mcu[3][0] * -32'h060) >> 8) + ((mcu[3][1] * -32'h051) >> 8) + ((mcu[3][2] * -32'h036) >> 8) + ((mcu[3][3] * -32'h013) >> 8) + ((mcu[3][4] * 32'h013) >> 8) + ((mcu[3][5] * 32'h036) >> 8) + ((mcu[3][6] * 32'h051) >> 8) + ((mcu[3][7] * 32'h060) >> 8) + ((mcu[4][0] * -32'h060) >> 8) + ((mcu[4][1] * -32'h051) >> 8) + ((mcu[4][2] * -32'h036) >> 8) + ((mcu[4][3] * -32'h013) >> 8) + ((mcu[4][4] * 32'h013) >> 8) + ((mcu[4][5] * 32'h036) >> 8) + ((mcu[4][6] * 32'h051) >> 8) + ((mcu[4][7] * 32'h060) >> 8) + ((mcu[5][0] * 32'h0e7) >> 8) + ((mcu[5][1] * 32'h0c4) >> 8) + ((mcu[5][2] * 32'h083) >> 8) + ((mcu[5][3] * 32'h02e) >> 8) + ((mcu[5][4] * -32'h02e) >> 8) + ((mcu[5][5] * -32'h083) >> 8) + ((mcu[5][6] * -32'h0c4) >> 8) + ((mcu[5][7] * -32'h0e7) >> 8) + ((mcu[6][0] * -32'h0e7) >> 8) + ((mcu[6][1] * -32'h0c4) >> 8) + ((mcu[6][2] * -32'h083) >> 8) + ((mcu[6][3] * -32'h02e) >> 8) + ((mcu[6][4] * 32'h02e) >> 8) + ((mcu[6][5] * 32'h083) >> 8) + ((mcu[6][6] * 32'h0c4) >> 8) + ((mcu[6][7] * 32'h0e7) >> 8) + ((mcu[7][0] * 32'h060) >> 8) + ((mcu[7][1] * 32'h051) >> 8) + ((mcu[7][2] * 32'h036) >> 8) + ((mcu[7][3] * 32'h013) >> 8) + ((mcu[7][4] * -32'h013) >> 8) + ((mcu[7][5] * -32'h036) >> 8) + ((mcu[7][6] * -32'h051) >> 8) + ((mcu[7][7] * -32'h060) >> 8);
	wire[63:0] cos62_term = ((mcu[0][0] * 32'h05a) >> 8) + ((mcu[0][1] * 32'h025) >> 8) + ((mcu[0][2] * -32'h025) >> 8) + ((mcu[0][3] * -32'h05a) >> 8) + ((mcu[0][4] * -32'h05a) >> 8) + ((mcu[0][5] * -32'h025) >> 8) + ((mcu[0][6] * 32'h025) >> 8) + ((mcu[0][7] * 32'h05a) >> 8) + ((mcu[1][0] * -32'h0da) >> 8) + ((mcu[1][1] * -32'h05a) >> 8) + ((mcu[1][2] * 32'h05a) >> 8) + ((mcu[1][3] * 32'h0da) >> 8) + ((mcu[1][4] * 32'h0da) >> 8) + ((mcu[1][5] * 32'h05a) >> 8) + ((mcu[1][6] * -32'h05a) >> 8) + ((mcu[1][7] * -32'h0da) >> 8) + ((mcu[2][0] * 32'h0da) >> 8) + ((mcu[2][1] * 32'h05a) >> 8) + ((mcu[2][2] * -32'h05a) >> 8) + ((mcu[2][3] * -32'h0da) >> 8) + ((mcu[2][4] * -32'h0da) >> 8) + ((mcu[2][5] * -32'h05a) >> 8) + ((mcu[2][6] * 32'h05a) >> 8) + ((mcu[2][7] * 32'h0da) >> 8) + ((mcu[3][0] * -32'h05a) >> 8) + ((mcu[3][1] * -32'h025) >> 8) + ((mcu[3][2] * 32'h025) >> 8) + ((mcu[3][3] * 32'h05a) >> 8) + ((mcu[3][4] * 32'h05a) >> 8) + ((mcu[3][5] * 32'h025) >> 8) + ((mcu[3][6] * -32'h025) >> 8) + ((mcu[3][7] * -32'h05a) >> 8) + ((mcu[4][0] * -32'h05a) >> 8) + ((mcu[4][1] * -32'h025) >> 8) + ((mcu[4][2] * 32'h025) >> 8) + ((mcu[4][3] * 32'h05a) >> 8) + ((mcu[4][4] * 32'h05a) >> 8) + ((mcu[4][5] * 32'h025) >> 8) + ((mcu[4][6] * -32'h025) >> 8) + ((mcu[4][7] * -32'h05a) >> 8) + ((mcu[5][0] * 32'h0da) >> 8) + ((mcu[5][1] * 32'h05a) >> 8) + ((mcu[5][2] * -32'h05a) >> 8) + ((mcu[5][3] * -32'h0da) >> 8) + ((mcu[5][4] * -32'h0da) >> 8) + ((mcu[5][5] * -32'h05a) >> 8) + ((mcu[5][6] * 32'h05a) >> 8) + ((mcu[5][7] * 32'h0da) >> 8) + ((mcu[6][0] * -32'h0da) >> 8) + ((mcu[6][1] * -32'h05a) >> 8) + ((mcu[6][2] * 32'h05a) >> 8) + ((mcu[6][3] * 32'h0da) >> 8) + ((mcu[6][4] * 32'h0da) >> 8) + ((mcu[6][5] * 32'h05a) >> 8) + ((mcu[6][6] * -32'h05a) >> 8) + ((mcu[6][7] * -32'h0da) >> 8) + ((mcu[7][0] * 32'h05a) >> 8) + ((mcu[7][1] * 32'h025) >> 8) + ((mcu[7][2] * -32'h025) >> 8) + ((mcu[7][3] * -32'h05a) >> 8) + ((mcu[7][4] * -32'h05a) >> 8) + ((mcu[7][5] * -32'h025) >> 8) + ((mcu[7][6] * 32'h025) >> 8) + ((mcu[7][7] * 32'h05a) >> 8);
	wire[63:0] cos63_term = ((mcu[0][0] * 32'h051) >> 8) + ((mcu[0][1] * -32'h013) >> 8) + ((mcu[0][2] * -32'h060) >> 8) + ((mcu[0][3] * -32'h036) >> 8) + ((mcu[0][4] * 32'h036) >> 8) + ((mcu[0][5] * 32'h060) >> 8) + ((mcu[0][6] * 32'h013) >> 8) + ((mcu[0][7] * -32'h051) >> 8) + ((mcu[1][0] * -32'h0c4) >> 8) + ((mcu[1][1] * 32'h02e) >> 8) + ((mcu[1][2] * 32'h0e7) >> 8) + ((mcu[1][3] * 32'h083) >> 8) + ((mcu[1][4] * -32'h083) >> 8) + ((mcu[1][5] * -32'h0e7) >> 8) + ((mcu[1][6] * -32'h02e) >> 8) + ((mcu[1][7] * 32'h0c4) >> 8) + ((mcu[2][0] * 32'h0c4) >> 8) + ((mcu[2][1] * -32'h02e) >> 8) + ((mcu[2][2] * -32'h0e7) >> 8) + ((mcu[2][3] * -32'h083) >> 8) + ((mcu[2][4] * 32'h083) >> 8) + ((mcu[2][5] * 32'h0e7) >> 8) + ((mcu[2][6] * 32'h02e) >> 8) + ((mcu[2][7] * -32'h0c4) >> 8) + ((mcu[3][0] * -32'h051) >> 8) + ((mcu[3][1] * 32'h013) >> 8) + ((mcu[3][2] * 32'h060) >> 8) + ((mcu[3][3] * 32'h036) >> 8) + ((mcu[3][4] * -32'h036) >> 8) + ((mcu[3][5] * -32'h060) >> 8) + ((mcu[3][6] * -32'h013) >> 8) + ((mcu[3][7] * 32'h051) >> 8) + ((mcu[4][0] * -32'h051) >> 8) + ((mcu[4][1] * 32'h013) >> 8) + ((mcu[4][2] * 32'h060) >> 8) + ((mcu[4][3] * 32'h036) >> 8) + ((mcu[4][4] * -32'h036) >> 8) + ((mcu[4][5] * -32'h060) >> 8) + ((mcu[4][6] * -32'h013) >> 8) + ((mcu[4][7] * 32'h051) >> 8) + ((mcu[5][0] * 32'h0c4) >> 8) + ((mcu[5][1] * -32'h02e) >> 8) + ((mcu[5][2] * -32'h0e7) >> 8) + ((mcu[5][3] * -32'h083) >> 8) + ((mcu[5][4] * 32'h083) >> 8) + ((mcu[5][5] * 32'h0e7) >> 8) + ((mcu[5][6] * 32'h02e) >> 8) + ((mcu[5][7] * -32'h0c4) >> 8) + ((mcu[6][0] * -32'h0c4) >> 8) + ((mcu[6][1] * 32'h02e) >> 8) + ((mcu[6][2] * 32'h0e7) >> 8) + ((mcu[6][3] * 32'h083) >> 8) + ((mcu[6][4] * -32'h083) >> 8) + ((mcu[6][5] * -32'h0e7) >> 8) + ((mcu[6][6] * -32'h02e) >> 8) + ((mcu[6][7] * 32'h0c4) >> 8) + ((mcu[7][0] * 32'h051) >> 8) + ((mcu[7][1] * -32'h013) >> 8) + ((mcu[7][2] * -32'h060) >> 8) + ((mcu[7][3] * -32'h036) >> 8) + ((mcu[7][4] * 32'h036) >> 8) + ((mcu[7][5] * 32'h060) >> 8) + ((mcu[7][6] * 32'h013) >> 8) + ((mcu[7][7] * -32'h051) >> 8);
	wire[63:0] cos64_term = ((mcu[0][0] * 32'h045) >> 8) + ((mcu[0][1] * -32'h045) >> 8) + ((mcu[0][2] * -32'h045) >> 8) + ((mcu[0][3] * 32'h045) >> 8) + ((mcu[0][4] * 32'h045) >> 8) + ((mcu[0][5] * -32'h045) >> 8) + ((mcu[0][6] * -32'h045) >> 8) + ((mcu[0][7] * 32'h045) >> 8) + ((mcu[1][0] * -32'h0a7) >> 8) + ((mcu[1][1] * 32'h0a7) >> 8) + ((mcu[1][2] * 32'h0a7) >> 8) + ((mcu[1][3] * -32'h0a7) >> 8) + ((mcu[1][4] * -32'h0a7) >> 8) + ((mcu[1][5] * 32'h0a7) >> 8) + ((mcu[1][6] * 32'h0a7) >> 8) + ((mcu[1][7] * -32'h0a7) >> 8) + ((mcu[2][0] * 32'h0a7) >> 8) + ((mcu[2][1] * -32'h0a7) >> 8) + ((mcu[2][2] * -32'h0a7) >> 8) + ((mcu[2][3] * 32'h0a7) >> 8) + ((mcu[2][4] * 32'h0a7) >> 8) + ((mcu[2][5] * -32'h0a7) >> 8) + ((mcu[2][6] * -32'h0a7) >> 8) + ((mcu[2][7] * 32'h0a7) >> 8) + ((mcu[3][0] * -32'h045) >> 8) + ((mcu[3][1] * 32'h045) >> 8) + ((mcu[3][2] * 32'h045) >> 8) + ((mcu[3][3] * -32'h045) >> 8) + ((mcu[3][4] * -32'h045) >> 8) + ((mcu[3][5] * 32'h045) >> 8) + ((mcu[3][6] * 32'h045) >> 8) + ((mcu[3][7] * -32'h045) >> 8) + ((mcu[4][0] * -32'h045) >> 8) + ((mcu[4][1] * 32'h045) >> 8) + ((mcu[4][2] * 32'h045) >> 8) + ((mcu[4][3] * -32'h045) >> 8) + ((mcu[4][4] * -32'h045) >> 8) + ((mcu[4][5] * 32'h045) >> 8) + ((mcu[4][6] * 32'h045) >> 8) + ((mcu[4][7] * -32'h045) >> 8) + ((mcu[5][0] * 32'h0a7) >> 8) + ((mcu[5][1] * -32'h0a7) >> 8) + ((mcu[5][2] * -32'h0a7) >> 8) + ((mcu[5][3] * 32'h0a7) >> 8) + ((mcu[5][4] * 32'h0a7) >> 8) + ((mcu[5][5] * -32'h0a7) >> 8) + ((mcu[5][6] * -32'h0a7) >> 8) + ((mcu[5][7] * 32'h0a7) >> 8) + ((mcu[6][0] * -32'h0a7) >> 8) + ((mcu[6][1] * 32'h0a7) >> 8) + ((mcu[6][2] * 32'h0a7) >> 8) + ((mcu[6][3] * -32'h0a7) >> 8) + ((mcu[6][4] * -32'h0a7) >> 8) + ((mcu[6][5] * 32'h0a7) >> 8) + ((mcu[6][6] * 32'h0a7) >> 8) + ((mcu[6][7] * -32'h0a7) >> 8) + ((mcu[7][0] * 32'h045) >> 8) + ((mcu[7][1] * -32'h045) >> 8) + ((mcu[7][2] * -32'h045) >> 8) + ((mcu[7][3] * 32'h045) >> 8) + ((mcu[7][4] * 32'h045) >> 8) + ((mcu[7][5] * -32'h045) >> 8) + ((mcu[7][6] * -32'h045) >> 8) + ((mcu[7][7] * 32'h045) >> 8);
	wire[63:0] cos65_term = ((mcu[0][0] * 32'h036) >> 8) + ((mcu[0][1] * -32'h060) >> 8) + ((mcu[0][2] * 32'h013) >> 8) + ((mcu[0][3] * 32'h051) >> 8) + ((mcu[0][4] * -32'h051) >> 8) + ((mcu[0][5] * -32'h013) >> 8) + ((mcu[0][6] * 32'h060) >> 8) + ((mcu[0][7] * -32'h036) >> 8) + ((mcu[1][0] * -32'h083) >> 8) + ((mcu[1][1] * 32'h0e7) >> 8) + ((mcu[1][2] * -32'h02e) >> 8) + ((mcu[1][3] * -32'h0c4) >> 8) + ((mcu[1][4] * 32'h0c4) >> 8) + ((mcu[1][5] * 32'h02e) >> 8) + ((mcu[1][6] * -32'h0e7) >> 8) + ((mcu[1][7] * 32'h083) >> 8) + ((mcu[2][0] * 32'h083) >> 8) + ((mcu[2][1] * -32'h0e7) >> 8) + ((mcu[2][2] * 32'h02e) >> 8) + ((mcu[2][3] * 32'h0c4) >> 8) + ((mcu[2][4] * -32'h0c4) >> 8) + ((mcu[2][5] * -32'h02e) >> 8) + ((mcu[2][6] * 32'h0e7) >> 8) + ((mcu[2][7] * -32'h083) >> 8) + ((mcu[3][0] * -32'h036) >> 8) + ((mcu[3][1] * 32'h060) >> 8) + ((mcu[3][2] * -32'h013) >> 8) + ((mcu[3][3] * -32'h051) >> 8) + ((mcu[3][4] * 32'h051) >> 8) + ((mcu[3][5] * 32'h013) >> 8) + ((mcu[3][6] * -32'h060) >> 8) + ((mcu[3][7] * 32'h036) >> 8) + ((mcu[4][0] * -32'h036) >> 8) + ((mcu[4][1] * 32'h060) >> 8) + ((mcu[4][2] * -32'h013) >> 8) + ((mcu[4][3] * -32'h051) >> 8) + ((mcu[4][4] * 32'h051) >> 8) + ((mcu[4][5] * 32'h013) >> 8) + ((mcu[4][6] * -32'h060) >> 8) + ((mcu[4][7] * 32'h036) >> 8) + ((mcu[5][0] * 32'h083) >> 8) + ((mcu[5][1] * -32'h0e7) >> 8) + ((mcu[5][2] * 32'h02e) >> 8) + ((mcu[5][3] * 32'h0c4) >> 8) + ((mcu[5][4] * -32'h0c4) >> 8) + ((mcu[5][5] * -32'h02e) >> 8) + ((mcu[5][6] * 32'h0e7) >> 8) + ((mcu[5][7] * -32'h083) >> 8) + ((mcu[6][0] * -32'h083) >> 8) + ((mcu[6][1] * 32'h0e7) >> 8) + ((mcu[6][2] * -32'h02e) >> 8) + ((mcu[6][3] * -32'h0c4) >> 8) + ((mcu[6][4] * 32'h0c4) >> 8) + ((mcu[6][5] * 32'h02e) >> 8) + ((mcu[6][6] * -32'h0e7) >> 8) + ((mcu[6][7] * 32'h083) >> 8) + ((mcu[7][0] * 32'h036) >> 8) + ((mcu[7][1] * -32'h060) >> 8) + ((mcu[7][2] * 32'h013) >> 8) + ((mcu[7][3] * 32'h051) >> 8) + ((mcu[7][4] * -32'h051) >> 8) + ((mcu[7][5] * -32'h013) >> 8) + ((mcu[7][6] * 32'h060) >> 8) + ((mcu[7][7] * -32'h036) >> 8);
	wire[63:0] cos66_term = ((mcu[0][0] * 32'h025) >> 8) + ((mcu[0][1] * -32'h05a) >> 8) + ((mcu[0][2] * 32'h05a) >> 8) + ((mcu[0][3] * -32'h025) >> 8) + ((mcu[0][4] * -32'h025) >> 8) + ((mcu[0][5] * 32'h05a) >> 8) + ((mcu[0][6] * -32'h05a) >> 8) + ((mcu[0][7] * 32'h025) >> 8) + ((mcu[1][0] * -32'h05a) >> 8) + ((mcu[1][1] * 32'h0da) >> 8) + ((mcu[1][2] * -32'h0da) >> 8) + ((mcu[1][3] * 32'h05a) >> 8) + ((mcu[1][4] * 32'h05a) >> 8) + ((mcu[1][5] * -32'h0da) >> 8) + ((mcu[1][6] * 32'h0da) >> 8) + ((mcu[1][7] * -32'h05a) >> 8) + ((mcu[2][0] * 32'h05a) >> 8) + ((mcu[2][1] * -32'h0da) >> 8) + ((mcu[2][2] * 32'h0da) >> 8) + ((mcu[2][3] * -32'h05a) >> 8) + ((mcu[2][4] * -32'h05a) >> 8) + ((mcu[2][5] * 32'h0da) >> 8) + ((mcu[2][6] * -32'h0da) >> 8) + ((mcu[2][7] * 32'h05a) >> 8) + ((mcu[3][0] * -32'h025) >> 8) + ((mcu[3][1] * 32'h05a) >> 8) + ((mcu[3][2] * -32'h05a) >> 8) + ((mcu[3][3] * 32'h025) >> 8) + ((mcu[3][4] * 32'h025) >> 8) + ((mcu[3][5] * -32'h05a) >> 8) + ((mcu[3][6] * 32'h05a) >> 8) + ((mcu[3][7] * -32'h025) >> 8) + ((mcu[4][0] * -32'h025) >> 8) + ((mcu[4][1] * 32'h05a) >> 8) + ((mcu[4][2] * -32'h05a) >> 8) + ((mcu[4][3] * 32'h025) >> 8) + ((mcu[4][4] * 32'h025) >> 8) + ((mcu[4][5] * -32'h05a) >> 8) + ((mcu[4][6] * 32'h05a) >> 8) + ((mcu[4][7] * -32'h025) >> 8) + ((mcu[5][0] * 32'h05a) >> 8) + ((mcu[5][1] * -32'h0da) >> 8) + ((mcu[5][2] * 32'h0da) >> 8) + ((mcu[5][3] * -32'h05a) >> 8) + ((mcu[5][4] * -32'h05a) >> 8) + ((mcu[5][5] * 32'h0da) >> 8) + ((mcu[5][6] * -32'h0da) >> 8) + ((mcu[5][7] * 32'h05a) >> 8) + ((mcu[6][0] * -32'h05a) >> 8) + ((mcu[6][1] * 32'h0da) >> 8) + ((mcu[6][2] * -32'h0da) >> 8) + ((mcu[6][3] * 32'h05a) >> 8) + ((mcu[6][4] * 32'h05a) >> 8) + ((mcu[6][5] * -32'h0da) >> 8) + ((mcu[6][6] * 32'h0da) >> 8) + ((mcu[6][7] * -32'h05a) >> 8) + ((mcu[7][0] * 32'h025) >> 8) + ((mcu[7][1] * -32'h05a) >> 8) + ((mcu[7][2] * 32'h05a) >> 8) + ((mcu[7][3] * -32'h025) >> 8) + ((mcu[7][4] * -32'h025) >> 8) + ((mcu[7][5] * 32'h05a) >> 8) + ((mcu[7][6] * -32'h05a) >> 8) + ((mcu[7][7] * 32'h025) >> 8);
	wire[63:0] cos67_term = ((mcu[0][0] * 32'h013) >> 8) + ((mcu[0][1] * -32'h036) >> 8) + ((mcu[0][2] * 32'h051) >> 8) + ((mcu[0][3] * -32'h060) >> 8) + ((mcu[0][4] * 32'h060) >> 8) + ((mcu[0][5] * -32'h051) >> 8) + ((mcu[0][6] * 32'h036) >> 8) + ((mcu[0][7] * -32'h013) >> 8) + ((mcu[1][0] * -32'h02e) >> 8) + ((mcu[1][1] * 32'h083) >> 8) + ((mcu[1][2] * -32'h0c4) >> 8) + ((mcu[1][3] * 32'h0e7) >> 8) + ((mcu[1][4] * -32'h0e7) >> 8) + ((mcu[1][5] * 32'h0c4) >> 8) + ((mcu[1][6] * -32'h083) >> 8) + ((mcu[1][7] * 32'h02e) >> 8) + ((mcu[2][0] * 32'h02e) >> 8) + ((mcu[2][1] * -32'h083) >> 8) + ((mcu[2][2] * 32'h0c4) >> 8) + ((mcu[2][3] * -32'h0e7) >> 8) + ((mcu[2][4] * 32'h0e7) >> 8) + ((mcu[2][5] * -32'h0c4) >> 8) + ((mcu[2][6] * 32'h083) >> 8) + ((mcu[2][7] * -32'h02e) >> 8) + ((mcu[3][0] * -32'h013) >> 8) + ((mcu[3][1] * 32'h036) >> 8) + ((mcu[3][2] * -32'h051) >> 8) + ((mcu[3][3] * 32'h060) >> 8) + ((mcu[3][4] * -32'h060) >> 8) + ((mcu[3][5] * 32'h051) >> 8) + ((mcu[3][6] * -32'h036) >> 8) + ((mcu[3][7] * 32'h013) >> 8) + ((mcu[4][0] * -32'h013) >> 8) + ((mcu[4][1] * 32'h036) >> 8) + ((mcu[4][2] * -32'h051) >> 8) + ((mcu[4][3] * 32'h060) >> 8) + ((mcu[4][4] * -32'h060) >> 8) + ((mcu[4][5] * 32'h051) >> 8) + ((mcu[4][6] * -32'h036) >> 8) + ((mcu[4][7] * 32'h013) >> 8) + ((mcu[5][0] * 32'h02e) >> 8) + ((mcu[5][1] * -32'h083) >> 8) + ((mcu[5][2] * 32'h0c4) >> 8) + ((mcu[5][3] * -32'h0e7) >> 8) + ((mcu[5][4] * 32'h0e7) >> 8) + ((mcu[5][5] * -32'h0c4) >> 8) + ((mcu[5][6] * 32'h083) >> 8) + ((mcu[5][7] * -32'h02e) >> 8) + ((mcu[6][0] * -32'h02e) >> 8) + ((mcu[6][1] * 32'h083) >> 8) + ((mcu[6][2] * -32'h0c4) >> 8) + ((mcu[6][3] * 32'h0e7) >> 8) + ((mcu[6][4] * -32'h0e7) >> 8) + ((mcu[6][5] * 32'h0c4) >> 8) + ((mcu[6][6] * -32'h083) >> 8) + ((mcu[6][7] * 32'h02e) >> 8) + ((mcu[7][0] * 32'h013) >> 8) + ((mcu[7][1] * -32'h036) >> 8) + ((mcu[7][2] * 32'h051) >> 8) + ((mcu[7][3] * -32'h060) >> 8) + ((mcu[7][4] * 32'h060) >> 8) + ((mcu[7][5] * -32'h051) >> 8) + ((mcu[7][6] * 32'h036) >> 8) + ((mcu[7][7] * -32'h013) >> 8);
	wire[63:0] cos70_term = ((mcu[0][0] * 32'h031) >> 8) + ((mcu[0][1] * 32'h031) >> 8) + ((mcu[0][2] * 32'h031) >> 8) + ((mcu[0][3] * 32'h031) >> 8) + ((mcu[0][4] * 32'h031) >> 8) + ((mcu[0][5] * 32'h031) >> 8) + ((mcu[0][6] * 32'h031) >> 8) + ((mcu[0][7] * 32'h031) >> 8) + ((mcu[1][0] * -32'h08e) >> 8) + ((mcu[1][1] * -32'h08e) >> 8) + ((mcu[1][2] * -32'h08e) >> 8) + ((mcu[1][3] * -32'h08e) >> 8) + ((mcu[1][4] * -32'h08e) >> 8) + ((mcu[1][5] * -32'h08e) >> 8) + ((mcu[1][6] * -32'h08e) >> 8) + ((mcu[1][7] * -32'h08e) >> 8) + ((mcu[2][0] * 32'h0d4) >> 8) + ((mcu[2][1] * 32'h0d4) >> 8) + ((mcu[2][2] * 32'h0d4) >> 8) + ((mcu[2][3] * 32'h0d4) >> 8) + ((mcu[2][4] * 32'h0d4) >> 8) + ((mcu[2][5] * 32'h0d4) >> 8) + ((mcu[2][6] * 32'h0d4) >> 8) + ((mcu[2][7] * 32'h0d4) >> 8) + ((mcu[3][0] * -32'h0fb) >> 8) + ((mcu[3][1] * -32'h0fb) >> 8) + ((mcu[3][2] * -32'h0fb) >> 8) + ((mcu[3][3] * -32'h0fb) >> 8) + ((mcu[3][4] * -32'h0fb) >> 8) + ((mcu[3][5] * -32'h0fb) >> 8) + ((mcu[3][6] * -32'h0fb) >> 8) + ((mcu[3][7] * -32'h0fb) >> 8) + ((mcu[4][0] * 32'h0fb) >> 8) + ((mcu[4][1] * 32'h0fb) >> 8) + ((mcu[4][2] * 32'h0fb) >> 8) + ((mcu[4][3] * 32'h0fb) >> 8) + ((mcu[4][4] * 32'h0fb) >> 8) + ((mcu[4][5] * 32'h0fb) >> 8) + ((mcu[4][6] * 32'h0fb) >> 8) + ((mcu[4][7] * 32'h0fb) >> 8) + ((mcu[5][0] * -32'h0d4) >> 8) + ((mcu[5][1] * -32'h0d4) >> 8) + ((mcu[5][2] * -32'h0d4) >> 8) + ((mcu[5][3] * -32'h0d4) >> 8) + ((mcu[5][4] * -32'h0d4) >> 8) + ((mcu[5][5] * -32'h0d4) >> 8) + ((mcu[5][6] * -32'h0d4) >> 8) + ((mcu[5][7] * -32'h0d4) >> 8) + ((mcu[6][0] * 32'h08e) >> 8) + ((mcu[6][1] * 32'h08e) >> 8) + ((mcu[6][2] * 32'h08e) >> 8) + ((mcu[6][3] * 32'h08e) >> 8) + ((mcu[6][4] * 32'h08e) >> 8) + ((mcu[6][5] * 32'h08e) >> 8) + ((mcu[6][6] * 32'h08e) >> 8) + ((mcu[6][7] * 32'h08e) >> 8) + ((mcu[7][0] * -32'h031) >> 8) + ((mcu[7][1] * -32'h031) >> 8) + ((mcu[7][2] * -32'h031) >> 8) + ((mcu[7][3] * -32'h031) >> 8) + ((mcu[7][4] * -32'h031) >> 8) + ((mcu[7][5] * -32'h031) >> 8) + ((mcu[7][6] * -32'h031) >> 8) + ((mcu[7][7] * -32'h031) >> 8);
	wire[63:0] cos71_term = ((mcu[0][0] * 32'h030) >> 8) + ((mcu[0][1] * 32'h029) >> 8) + ((mcu[0][2] * 32'h01b) >> 8) + ((mcu[0][3] * 32'h009) >> 8) + ((mcu[0][4] * -32'h009) >> 8) + ((mcu[0][5] * -32'h01b) >> 8) + ((mcu[0][6] * -32'h029) >> 8) + ((mcu[0][7] * -32'h030) >> 8) + ((mcu[1][0] * -32'h08b) >> 8) + ((mcu[1][1] * -32'h076) >> 8) + ((mcu[1][2] * -32'h04f) >> 8) + ((mcu[1][3] * -32'h01b) >> 8) + ((mcu[1][4] * 32'h01b) >> 8) + ((mcu[1][5] * 32'h04f) >> 8) + ((mcu[1][6] * 32'h076) >> 8) + ((mcu[1][7] * 32'h08b) >> 8) + ((mcu[2][0] * 32'h0d0) >> 8) + ((mcu[2][1] * 32'h0b0) >> 8) + ((mcu[2][2] * 32'h076) >> 8) + ((mcu[2][3] * 32'h029) >> 8) + ((mcu[2][4] * -32'h029) >> 8) + ((mcu[2][5] * -32'h076) >> 8) + ((mcu[2][6] * -32'h0b0) >> 8) + ((mcu[2][7] * -32'h0d0) >> 8) + ((mcu[3][0] * -32'h0f6) >> 8) + ((mcu[3][1] * -32'h0d0) >> 8) + ((mcu[3][2] * -32'h08b) >> 8) + ((mcu[3][3] * -32'h030) >> 8) + ((mcu[3][4] * 32'h030) >> 8) + ((mcu[3][5] * 32'h08b) >> 8) + ((mcu[3][6] * 32'h0d0) >> 8) + ((mcu[3][7] * 32'h0f6) >> 8) + ((mcu[4][0] * 32'h0f6) >> 8) + ((mcu[4][1] * 32'h0d0) >> 8) + ((mcu[4][2] * 32'h08b) >> 8) + ((mcu[4][3] * 32'h030) >> 8) + ((mcu[4][4] * -32'h030) >> 8) + ((mcu[4][5] * -32'h08b) >> 8) + ((mcu[4][6] * -32'h0d0) >> 8) + ((mcu[4][7] * -32'h0f6) >> 8) + ((mcu[5][0] * -32'h0d0) >> 8) + ((mcu[5][1] * -32'h0b0) >> 8) + ((mcu[5][2] * -32'h076) >> 8) + ((mcu[5][3] * -32'h029) >> 8) + ((mcu[5][4] * 32'h029) >> 8) + ((mcu[5][5] * 32'h076) >> 8) + ((mcu[5][6] * 32'h0b0) >> 8) + ((mcu[5][7] * 32'h0d0) >> 8) + ((mcu[6][0] * 32'h08b) >> 8) + ((mcu[6][1] * 32'h076) >> 8) + ((mcu[6][2] * 32'h04f) >> 8) + ((mcu[6][3] * 32'h01b) >> 8) + ((mcu[6][4] * -32'h01b) >> 8) + ((mcu[6][5] * -32'h04f) >> 8) + ((mcu[6][6] * -32'h076) >> 8) + ((mcu[6][7] * -32'h08b) >> 8) + ((mcu[7][0] * -32'h030) >> 8) + ((mcu[7][1] * -32'h029) >> 8) + ((mcu[7][2] * -32'h01b) >> 8) + ((mcu[7][3] * -32'h009) >> 8) + ((mcu[7][4] * 32'h009) >> 8) + ((mcu[7][5] * 32'h01b) >> 8) + ((mcu[7][6] * 32'h029) >> 8) + ((mcu[7][7] * 32'h030) >> 8);
	wire[63:0] cos72_term = ((mcu[0][0] * 32'h02e) >> 8) + ((mcu[0][1] * 32'h013) >> 8) + ((mcu[0][2] * -32'h013) >> 8) + ((mcu[0][3] * -32'h02e) >> 8) + ((mcu[0][4] * -32'h02e) >> 8) + ((mcu[0][5] * -32'h013) >> 8) + ((mcu[0][6] * 32'h013) >> 8) + ((mcu[0][7] * 32'h02e) >> 8) + ((mcu[1][0] * -32'h083) >> 8) + ((mcu[1][1] * -32'h036) >> 8) + ((mcu[1][2] * 32'h036) >> 8) + ((mcu[1][3] * 32'h083) >> 8) + ((mcu[1][4] * 32'h083) >> 8) + ((mcu[1][5] * 32'h036) >> 8) + ((mcu[1][6] * -32'h036) >> 8) + ((mcu[1][7] * -32'h083) >> 8) + ((mcu[2][0] * 32'h0c4) >> 8) + ((mcu[2][1] * 32'h051) >> 8) + ((mcu[2][2] * -32'h051) >> 8) + ((mcu[2][3] * -32'h0c4) >> 8) + ((mcu[2][4] * -32'h0c4) >> 8) + ((mcu[2][5] * -32'h051) >> 8) + ((mcu[2][6] * 32'h051) >> 8) + ((mcu[2][7] * 32'h0c4) >> 8) + ((mcu[3][0] * -32'h0e7) >> 8) + ((mcu[3][1] * -32'h060) >> 8) + ((mcu[3][2] * 32'h060) >> 8) + ((mcu[3][3] * 32'h0e7) >> 8) + ((mcu[3][4] * 32'h0e7) >> 8) + ((mcu[3][5] * 32'h060) >> 8) + ((mcu[3][6] * -32'h060) >> 8) + ((mcu[3][7] * -32'h0e7) >> 8) + ((mcu[4][0] * 32'h0e7) >> 8) + ((mcu[4][1] * 32'h060) >> 8) + ((mcu[4][2] * -32'h060) >> 8) + ((mcu[4][3] * -32'h0e7) >> 8) + ((mcu[4][4] * -32'h0e7) >> 8) + ((mcu[4][5] * -32'h060) >> 8) + ((mcu[4][6] * 32'h060) >> 8) + ((mcu[4][7] * 32'h0e7) >> 8) + ((mcu[5][0] * -32'h0c4) >> 8) + ((mcu[5][1] * -32'h051) >> 8) + ((mcu[5][2] * 32'h051) >> 8) + ((mcu[5][3] * 32'h0c4) >> 8) + ((mcu[5][4] * 32'h0c4) >> 8) + ((mcu[5][5] * 32'h051) >> 8) + ((mcu[5][6] * -32'h051) >> 8) + ((mcu[5][7] * -32'h0c4) >> 8) + ((mcu[6][0] * 32'h083) >> 8) + ((mcu[6][1] * 32'h036) >> 8) + ((mcu[6][2] * -32'h036) >> 8) + ((mcu[6][3] * -32'h083) >> 8) + ((mcu[6][4] * -32'h083) >> 8) + ((mcu[6][5] * -32'h036) >> 8) + ((mcu[6][6] * 32'h036) >> 8) + ((mcu[6][7] * 32'h083) >> 8) + ((mcu[7][0] * -32'h02e) >> 8) + ((mcu[7][1] * -32'h013) >> 8) + ((mcu[7][2] * 32'h013) >> 8) + ((mcu[7][3] * 32'h02e) >> 8) + ((mcu[7][4] * 32'h02e) >> 8) + ((mcu[7][5] * 32'h013) >> 8) + ((mcu[7][6] * -32'h013) >> 8) + ((mcu[7][7] * -32'h02e) >> 8);
	wire[63:0] cos73_term = ((mcu[0][0] * 32'h029) >> 8) + ((mcu[0][1] * -32'h009) >> 8) + ((mcu[0][2] * -32'h030) >> 8) + ((mcu[0][3] * -32'h01b) >> 8) + ((mcu[0][4] * 32'h01b) >> 8) + ((mcu[0][5] * 32'h030) >> 8) + ((mcu[0][6] * 32'h009) >> 8) + ((mcu[0][7] * -32'h029) >> 8) + ((mcu[1][0] * -32'h076) >> 8) + ((mcu[1][1] * 32'h01b) >> 8) + ((mcu[1][2] * 32'h08b) >> 8) + ((mcu[1][3] * 32'h04f) >> 8) + ((mcu[1][4] * -32'h04f) >> 8) + ((mcu[1][5] * -32'h08b) >> 8) + ((mcu[1][6] * -32'h01b) >> 8) + ((mcu[1][7] * 32'h076) >> 8) + ((mcu[2][0] * 32'h0b0) >> 8) + ((mcu[2][1] * -32'h029) >> 8) + ((mcu[2][2] * -32'h0d0) >> 8) + ((mcu[2][3] * -32'h076) >> 8) + ((mcu[2][4] * 32'h076) >> 8) + ((mcu[2][5] * 32'h0d0) >> 8) + ((mcu[2][6] * 32'h029) >> 8) + ((mcu[2][7] * -32'h0b0) >> 8) + ((mcu[3][0] * -32'h0d0) >> 8) + ((mcu[3][1] * 32'h030) >> 8) + ((mcu[3][2] * 32'h0f6) >> 8) + ((mcu[3][3] * 32'h08b) >> 8) + ((mcu[3][4] * -32'h08b) >> 8) + ((mcu[3][5] * -32'h0f6) >> 8) + ((mcu[3][6] * -32'h030) >> 8) + ((mcu[3][7] * 32'h0d0) >> 8) + ((mcu[4][0] * 32'h0d0) >> 8) + ((mcu[4][1] * -32'h030) >> 8) + ((mcu[4][2] * -32'h0f6) >> 8) + ((mcu[4][3] * -32'h08b) >> 8) + ((mcu[4][4] * 32'h08b) >> 8) + ((mcu[4][5] * 32'h0f6) >> 8) + ((mcu[4][6] * 32'h030) >> 8) + ((mcu[4][7] * -32'h0d0) >> 8) + ((mcu[5][0] * -32'h0b0) >> 8) + ((mcu[5][1] * 32'h029) >> 8) + ((mcu[5][2] * 32'h0d0) >> 8) + ((mcu[5][3] * 32'h076) >> 8) + ((mcu[5][4] * -32'h076) >> 8) + ((mcu[5][5] * -32'h0d0) >> 8) + ((mcu[5][6] * -32'h029) >> 8) + ((mcu[5][7] * 32'h0b0) >> 8) + ((mcu[6][0] * 32'h076) >> 8) + ((mcu[6][1] * -32'h01b) >> 8) + ((mcu[6][2] * -32'h08b) >> 8) + ((mcu[6][3] * -32'h04f) >> 8) + ((mcu[6][4] * 32'h04f) >> 8) + ((mcu[6][5] * 32'h08b) >> 8) + ((mcu[6][6] * 32'h01b) >> 8) + ((mcu[6][7] * -32'h076) >> 8) + ((mcu[7][0] * -32'h029) >> 8) + ((mcu[7][1] * 32'h009) >> 8) + ((mcu[7][2] * 32'h030) >> 8) + ((mcu[7][3] * 32'h01b) >> 8) + ((mcu[7][4] * -32'h01b) >> 8) + ((mcu[7][5] * -32'h030) >> 8) + ((mcu[7][6] * -32'h009) >> 8) + ((mcu[7][7] * 32'h029) >> 8);
	wire[63:0] cos74_term = ((mcu[0][0] * 32'h023) >> 8) + ((mcu[0][1] * -32'h023) >> 8) + ((mcu[0][2] * -32'h023) >> 8) + ((mcu[0][3] * 32'h023) >> 8) + ((mcu[0][4] * 32'h023) >> 8) + ((mcu[0][5] * -32'h023) >> 8) + ((mcu[0][6] * -32'h023) >> 8) + ((mcu[0][7] * 32'h023) >> 8) + ((mcu[1][0] * -32'h064) >> 8) + ((mcu[1][1] * 32'h064) >> 8) + ((mcu[1][2] * 32'h064) >> 8) + ((mcu[1][3] * -32'h064) >> 8) + ((mcu[1][4] * -32'h064) >> 8) + ((mcu[1][5] * 32'h064) >> 8) + ((mcu[1][6] * 32'h064) >> 8) + ((mcu[1][7] * -32'h064) >> 8) + ((mcu[2][0] * 32'h096) >> 8) + ((mcu[2][1] * -32'h096) >> 8) + ((mcu[2][2] * -32'h096) >> 8) + ((mcu[2][3] * 32'h096) >> 8) + ((mcu[2][4] * 32'h096) >> 8) + ((mcu[2][5] * -32'h096) >> 8) + ((mcu[2][6] * -32'h096) >> 8) + ((mcu[2][7] * 32'h096) >> 8) + ((mcu[3][0] * -32'h0b1) >> 8) + ((mcu[3][1] * 32'h0b1) >> 8) + ((mcu[3][2] * 32'h0b1) >> 8) + ((mcu[3][3] * -32'h0b1) >> 8) + ((mcu[3][4] * -32'h0b1) >> 8) + ((mcu[3][5] * 32'h0b1) >> 8) + ((mcu[3][6] * 32'h0b1) >> 8) + ((mcu[3][7] * -32'h0b1) >> 8) + ((mcu[4][0] * 32'h0b1) >> 8) + ((mcu[4][1] * -32'h0b1) >> 8) + ((mcu[4][2] * -32'h0b1) >> 8) + ((mcu[4][3] * 32'h0b1) >> 8) + ((mcu[4][4] * 32'h0b1) >> 8) + ((mcu[4][5] * -32'h0b1) >> 8) + ((mcu[4][6] * -32'h0b1) >> 8) + ((mcu[4][7] * 32'h0b1) >> 8) + ((mcu[5][0] * -32'h096) >> 8) + ((mcu[5][1] * 32'h096) >> 8) + ((mcu[5][2] * 32'h096) >> 8) + ((mcu[5][3] * -32'h096) >> 8) + ((mcu[5][4] * -32'h096) >> 8) + ((mcu[5][5] * 32'h096) >> 8) + ((mcu[5][6] * 32'h096) >> 8) + ((mcu[5][7] * -32'h096) >> 8) + ((mcu[6][0] * 32'h064) >> 8) + ((mcu[6][1] * -32'h064) >> 8) + ((mcu[6][2] * -32'h064) >> 8) + ((mcu[6][3] * 32'h064) >> 8) + ((mcu[6][4] * 32'h064) >> 8) + ((mcu[6][5] * -32'h064) >> 8) + ((mcu[6][6] * -32'h064) >> 8) + ((mcu[6][7] * 32'h064) >> 8) + ((mcu[7][0] * -32'h023) >> 8) + ((mcu[7][1] * 32'h023) >> 8) + ((mcu[7][2] * 32'h023) >> 8) + ((mcu[7][3] * -32'h023) >> 8) + ((mcu[7][4] * -32'h023) >> 8) + ((mcu[7][5] * 32'h023) >> 8) + ((mcu[7][6] * 32'h023) >> 8) + ((mcu[7][7] * -32'h023) >> 8);
	wire[63:0] cos75_term = ((mcu[0][0] * 32'h01b) >> 8) + ((mcu[0][1] * -32'h030) >> 8) + ((mcu[0][2] * 32'h009) >> 8) + ((mcu[0][3] * 32'h029) >> 8) + ((mcu[0][4] * -32'h029) >> 8) + ((mcu[0][5] * -32'h009) >> 8) + ((mcu[0][6] * 32'h030) >> 8) + ((mcu[0][7] * -32'h01b) >> 8) + ((mcu[1][0] * -32'h04f) >> 8) + ((mcu[1][1] * 32'h08b) >> 8) + ((mcu[1][2] * -32'h01b) >> 8) + ((mcu[1][3] * -32'h076) >> 8) + ((mcu[1][4] * 32'h076) >> 8) + ((mcu[1][5] * 32'h01b) >> 8) + ((mcu[1][6] * -32'h08b) >> 8) + ((mcu[1][7] * 32'h04f) >> 8) + ((mcu[2][0] * 32'h076) >> 8) + ((mcu[2][1] * -32'h0d0) >> 8) + ((mcu[2][2] * 32'h029) >> 8) + ((mcu[2][3] * 32'h0b0) >> 8) + ((mcu[2][4] * -32'h0b0) >> 8) + ((mcu[2][5] * -32'h029) >> 8) + ((mcu[2][6] * 32'h0d0) >> 8) + ((mcu[2][7] * -32'h076) >> 8) + ((mcu[3][0] * -32'h08b) >> 8) + ((mcu[3][1] * 32'h0f6) >> 8) + ((mcu[3][2] * -32'h030) >> 8) + ((mcu[3][3] * -32'h0d0) >> 8) + ((mcu[3][4] * 32'h0d0) >> 8) + ((mcu[3][5] * 32'h030) >> 8) + ((mcu[3][6] * -32'h0f6) >> 8) + ((mcu[3][7] * 32'h08b) >> 8) + ((mcu[4][0] * 32'h08b) >> 8) + ((mcu[4][1] * -32'h0f6) >> 8) + ((mcu[4][2] * 32'h030) >> 8) + ((mcu[4][3] * 32'h0d0) >> 8) + ((mcu[4][4] * -32'h0d0) >> 8) + ((mcu[4][5] * -32'h030) >> 8) + ((mcu[4][6] * 32'h0f6) >> 8) + ((mcu[4][7] * -32'h08b) >> 8) + ((mcu[5][0] * -32'h076) >> 8) + ((mcu[5][1] * 32'h0d0) >> 8) + ((mcu[5][2] * -32'h029) >> 8) + ((mcu[5][3] * -32'h0b0) >> 8) + ((mcu[5][4] * 32'h0b0) >> 8) + ((mcu[5][5] * 32'h029) >> 8) + ((mcu[5][6] * -32'h0d0) >> 8) + ((mcu[5][7] * 32'h076) >> 8) + ((mcu[6][0] * 32'h04f) >> 8) + ((mcu[6][1] * -32'h08b) >> 8) + ((mcu[6][2] * 32'h01b) >> 8) + ((mcu[6][3] * 32'h076) >> 8) + ((mcu[6][4] * -32'h076) >> 8) + ((mcu[6][5] * -32'h01b) >> 8) + ((mcu[6][6] * 32'h08b) >> 8) + ((mcu[6][7] * -32'h04f) >> 8) + ((mcu[7][0] * -32'h01b) >> 8) + ((mcu[7][1] * 32'h030) >> 8) + ((mcu[7][2] * -32'h009) >> 8) + ((mcu[7][3] * -32'h029) >> 8) + ((mcu[7][4] * 32'h029) >> 8) + ((mcu[7][5] * 32'h009) >> 8) + ((mcu[7][6] * -32'h030) >> 8) + ((mcu[7][7] * 32'h01b) >> 8);
	wire[63:0] cos76_term = ((mcu[0][0] * 32'h013) >> 8) + ((mcu[0][1] * -32'h02e) >> 8) + ((mcu[0][2] * 32'h02e) >> 8) + ((mcu[0][3] * -32'h013) >> 8) + ((mcu[0][4] * -32'h013) >> 8) + ((mcu[0][5] * 32'h02e) >> 8) + ((mcu[0][6] * -32'h02e) >> 8) + ((mcu[0][7] * 32'h013) >> 8) + ((mcu[1][0] * -32'h036) >> 8) + ((mcu[1][1] * 32'h083) >> 8) + ((mcu[1][2] * -32'h083) >> 8) + ((mcu[1][3] * 32'h036) >> 8) + ((mcu[1][4] * 32'h036) >> 8) + ((mcu[1][5] * -32'h083) >> 8) + ((mcu[1][6] * 32'h083) >> 8) + ((mcu[1][7] * -32'h036) >> 8) + ((mcu[2][0] * 32'h051) >> 8) + ((mcu[2][1] * -32'h0c4) >> 8) + ((mcu[2][2] * 32'h0c4) >> 8) + ((mcu[2][3] * -32'h051) >> 8) + ((mcu[2][4] * -32'h051) >> 8) + ((mcu[2][5] * 32'h0c4) >> 8) + ((mcu[2][6] * -32'h0c4) >> 8) + ((mcu[2][7] * 32'h051) >> 8) + ((mcu[3][0] * -32'h060) >> 8) + ((mcu[3][1] * 32'h0e7) >> 8) + ((mcu[3][2] * -32'h0e7) >> 8) + ((mcu[3][3] * 32'h060) >> 8) + ((mcu[3][4] * 32'h060) >> 8) + ((mcu[3][5] * -32'h0e7) >> 8) + ((mcu[3][6] * 32'h0e7) >> 8) + ((mcu[3][7] * -32'h060) >> 8) + ((mcu[4][0] * 32'h060) >> 8) + ((mcu[4][1] * -32'h0e7) >> 8) + ((mcu[4][2] * 32'h0e7) >> 8) + ((mcu[4][3] * -32'h060) >> 8) + ((mcu[4][4] * -32'h060) >> 8) + ((mcu[4][5] * 32'h0e7) >> 8) + ((mcu[4][6] * -32'h0e7) >> 8) + ((mcu[4][7] * 32'h060) >> 8) + ((mcu[5][0] * -32'h051) >> 8) + ((mcu[5][1] * 32'h0c4) >> 8) + ((mcu[5][2] * -32'h0c4) >> 8) + ((mcu[5][3] * 32'h051) >> 8) + ((mcu[5][4] * 32'h051) >> 8) + ((mcu[5][5] * -32'h0c4) >> 8) + ((mcu[5][6] * 32'h0c4) >> 8) + ((mcu[5][7] * -32'h051) >> 8) + ((mcu[6][0] * 32'h036) >> 8) + ((mcu[6][1] * -32'h083) >> 8) + ((mcu[6][2] * 32'h083) >> 8) + ((mcu[6][3] * -32'h036) >> 8) + ((mcu[6][4] * -32'h036) >> 8) + ((mcu[6][5] * 32'h083) >> 8) + ((mcu[6][6] * -32'h083) >> 8) + ((mcu[6][7] * 32'h036) >> 8) + ((mcu[7][0] * -32'h013) >> 8) + ((mcu[7][1] * 32'h02e) >> 8) + ((mcu[7][2] * -32'h02e) >> 8) + ((mcu[7][3] * 32'h013) >> 8) + ((mcu[7][4] * 32'h013) >> 8) + ((mcu[7][5] * -32'h02e) >> 8) + ((mcu[7][6] * 32'h02e) >> 8) + ((mcu[7][7] * -32'h013) >> 8);
	wire[63:0] cos77_term = ((mcu[0][0] * 32'h009) >> 8) + ((mcu[0][1] * -32'h01b) >> 8) + ((mcu[0][2] * 32'h029) >> 8) + ((mcu[0][3] * -32'h030) >> 8) + ((mcu[0][4] * 32'h030) >> 8) + ((mcu[0][5] * -32'h029) >> 8) + ((mcu[0][6] * 32'h01b) >> 8) + ((mcu[0][7] * -32'h009) >> 8) + ((mcu[1][0] * -32'h01b) >> 8) + ((mcu[1][1] * 32'h04f) >> 8) + ((mcu[1][2] * -32'h076) >> 8) + ((mcu[1][3] * 32'h08b) >> 8) + ((mcu[1][4] * -32'h08b) >> 8) + ((mcu[1][5] * 32'h076) >> 8) + ((mcu[1][6] * -32'h04f) >> 8) + ((mcu[1][7] * 32'h01b) >> 8) + ((mcu[2][0] * 32'h029) >> 8) + ((mcu[2][1] * -32'h076) >> 8) + ((mcu[2][2] * 32'h0b0) >> 8) + ((mcu[2][3] * -32'h0d0) >> 8) + ((mcu[2][4] * 32'h0d0) >> 8) + ((mcu[2][5] * -32'h0b0) >> 8) + ((mcu[2][6] * 32'h076) >> 8) + ((mcu[2][7] * -32'h029) >> 8) + ((mcu[3][0] * -32'h030) >> 8) + ((mcu[3][1] * 32'h08b) >> 8) + ((mcu[3][2] * -32'h0d0) >> 8) + ((mcu[3][3] * 32'h0f6) >> 8) + ((mcu[3][4] * -32'h0f6) >> 8) + ((mcu[3][5] * 32'h0d0) >> 8) + ((mcu[3][6] * -32'h08b) >> 8) + ((mcu[3][7] * 32'h030) >> 8) + ((mcu[4][0] * 32'h030) >> 8) + ((mcu[4][1] * -32'h08b) >> 8) + ((mcu[4][2] * 32'h0d0) >> 8) + ((mcu[4][3] * -32'h0f6) >> 8) + ((mcu[4][4] * 32'h0f6) >> 8) + ((mcu[4][5] * -32'h0d0) >> 8) + ((mcu[4][6] * 32'h08b) >> 8) + ((mcu[4][7] * -32'h030) >> 8) + ((mcu[5][0] * -32'h029) >> 8) + ((mcu[5][1] * 32'h076) >> 8) + ((mcu[5][2] * -32'h0b0) >> 8) + ((mcu[5][3] * 32'h0d0) >> 8) + ((mcu[5][4] * -32'h0d0) >> 8) + ((mcu[5][5] * 32'h0b0) >> 8) + ((mcu[5][6] * -32'h076) >> 8) + ((mcu[5][7] * 32'h029) >> 8) + ((mcu[6][0] * 32'h01b) >> 8) + ((mcu[6][1] * -32'h04f) >> 8) + ((mcu[6][2] * 32'h076) >> 8) + ((mcu[6][3] * -32'h08b) >> 8) + ((mcu[6][4] * 32'h08b) >> 8) + ((mcu[6][5] * -32'h076) >> 8) + ((mcu[6][6] * 32'h04f) >> 8) + ((mcu[6][7] * -32'h01b) >> 8) + ((mcu[7][0] * -32'h009) >> 8) + ((mcu[7][1] * 32'h01b) >> 8) + ((mcu[7][2] * -32'h029) >> 8) + ((mcu[7][3] * 32'h030) >> 8) + ((mcu[7][4] * -32'h030) >> 8) + ((mcu[7][5] * 32'h029) >> 8) + ((mcu[7][6] * -32'h01b) >> 8) + ((mcu[7][7] * 32'h009) >> 8);
	
	wire[63:0] cos00_term_quantized = (cos00_term[31:0] / 32'h10_00) << 8;
	wire[63:0] cos01_term_quantized = (cos01_term[31:0] / 32'h0B_00) << 8;
	wire[63:0] cos02_term_quantized = (cos02_term[31:0] / 32'h0A_00) << 8;
	wire[63:0] cos03_term_quantized = (cos03_term[31:0] / 32'h10_00) << 8;
	wire[63:0] cos04_term_quantized = (cos04_term[31:0] / 32'h18_00) << 8;
	wire[63:0] cos05_term_quantized = (cos05_term[31:0] / 32'h28_00) << 8;
	wire[63:0] cos06_term_quantized = (cos06_term[31:0] / 32'h33_00) << 8;
	wire[63:0] cos07_term_quantized = (cos07_term[31:0] / 32'h3d_00) << 8;
	wire[63:0] cos10_term_quantized = (cos10_term[31:0] / 32'h0c_00) << 8;
	wire[63:0] cos11_term_quantized = (cos11_term[31:0] / 32'h0c_00) << 8;
	wire[63:0] cos12_term_quantized = (cos12_term[31:0] / 32'h0e_00) << 8;
	wire[63:0] cos13_term_quantized = (cos13_term[31:0] / 32'h13_00) << 8;
	wire[63:0] cos14_term_quantized = (cos14_term[31:0] / 32'h1a_00) << 8;
	wire[63:0] cos15_term_quantized = (cos15_term[31:0] / 32'h3a_00) << 8;
	wire[63:0] cos16_term_quantized = (cos16_term[31:0] / 32'h3c_00) << 8;
	wire[63:0] cos17_term_quantized = (cos17_term[31:0] / 32'h37_00) << 8;
	wire[63:0] cos20_term_quantized = (cos20_term[31:0] / 32'h0e_00) << 8;
	wire[63:0] cos21_term_quantized = (cos21_term[31:0] / 32'h0d_00) << 8;
	wire[63:0] cos22_term_quantized = (cos22_term[31:0] / 32'h10_00) << 8;
	wire[63:0] cos23_term_quantized = (cos23_term[31:0] / 32'h18_00) << 8;
	wire[63:0] cos24_term_quantized = (cos24_term[31:0] / 32'h28_00) << 8;
	wire[63:0] cos25_term_quantized = (cos25_term[31:0] / 32'h39_00) << 8;
	wire[63:0] cos26_term_quantized = (cos26_term[31:0] / 32'h45_00) << 8;
	wire[63:0] cos27_term_quantized = (cos27_term[31:0] / 32'h38_00) << 8;
	wire[63:0] cos30_term_quantized = (cos30_term[31:0] / 32'h0e_00) << 8;
	wire[63:0] cos31_term_quantized = (cos31_term[31:0] / 32'h11_00) << 8;
	wire[63:0] cos32_term_quantized = (cos32_term[31:0] / 32'h16_00) << 8;
	wire[63:0] cos33_term_quantized = (cos33_term[31:0] / 32'h1d_00) << 8;
	wire[63:0] cos34_term_quantized = (cos34_term[31:0] / 32'h33_00) << 8;
	wire[63:0] cos35_term_quantized = (cos35_term[31:0] / 32'h57_00) << 8;
	wire[63:0] cos36_term_quantized = (cos36_term[31:0] / 32'h57_00) << 8;
	wire[63:0] cos37_term_quantized = (cos37_term[31:0] / 32'h3e_00) << 8;
	wire[63:0] cos40_term_quantized = (cos40_term[31:0] / 32'h12_00) << 8;
	wire[63:0] cos41_term_quantized = (cos41_term[31:0] / 32'h16_00) << 8;
	wire[63:0] cos42_term_quantized = (cos42_term[31:0] / 32'h25_00) << 8;
	wire[63:0] cos43_term_quantized = (cos43_term[31:0] / 32'h38_00) << 8;
	wire[63:0] cos44_term_quantized = (cos44_term[31:0] / 32'h44_00) << 8;
	wire[63:0] cos45_term_quantized = (cos45_term[31:0] / 32'h6d_00) << 8;
	wire[63:0] cos46_term_quantized = (cos46_term[31:0] / 32'h67_00) << 8;
	wire[63:0] cos47_term_quantized = (cos47_term[31:0] / 32'h4d_00) << 8;
	wire[63:0] cos50_term_quantized = (cos50_term[31:0] / 32'h18_00) << 8;
	wire[63:0] cos51_term_quantized = (cos51_term[31:0] / 32'h23_00) << 8;
	wire[63:0] cos52_term_quantized = (cos52_term[31:0] / 32'h37_00) << 8;
	wire[63:0] cos53_term_quantized = (cos53_term[31:0] / 32'h40_00) << 8;
	wire[63:0] cos54_term_quantized = (cos54_term[31:0] / 32'h51_00) << 8;
	wire[63:0] cos55_term_quantized = (cos55_term[31:0] / 32'h68_00) << 8;
	wire[63:0] cos56_term_quantized = (cos56_term[31:0] / 32'h71_00) << 8;
	wire[63:0] cos57_term_quantized = (cos57_term[31:0] / 32'h5c_00) << 8;
	wire[63:0] cos60_term_quantized = (cos60_term[31:0] / 32'h31_00) << 8;
	wire[63:0] cos61_term_quantized = (cos61_term[31:0] / 32'h40_00) << 8;
	wire[63:0] cos62_term_quantized = (cos62_term[31:0] / 32'h4e_00) << 8;
	wire[63:0] cos63_term_quantized = (cos63_term[31:0] / 32'h57_00) << 8;
	wire[63:0] cos64_term_quantized = (cos64_term[31:0] / 32'h67_00) << 8;
	wire[63:0] cos65_term_quantized = (cos65_term[31:0] / 32'h79_00) << 8;
	wire[63:0] cos66_term_quantized = (cos66_term[31:0] / 32'h78_00) << 8;
	wire[63:0] cos67_term_quantized = (cos67_term[31:0] / 32'h65_00) << 8;
	wire[63:0] cos70_term_quantized = (cos70_term[31:0] / 32'h48_00) << 8;
	wire[63:0] cos71_term_quantized = (cos71_term[31:0] / 32'h5c_00) << 8;
	wire[63:0] cos72_term_quantized = (cos72_term[31:0] / 32'h5f_00) << 8;
	wire[63:0] cos73_term_quantized = (cos73_term[31:0] / 32'h62_00) << 8;
	wire[63:0] cos74_term_quantized = (cos74_term[31:0] / 32'h70_00) << 8;
	wire[63:0] cos75_term_quantized = (cos75_term[31:0] / 32'h64_00) << 8;
	wire[63:0] cos76_term_quantized = (cos76_term[31:0] / 32'h67_00) << 8;
	wire[63:0] cos77_term_quantized = (cos77_term[31:0] / 32'h63_00) << 8;

	always_comb begin
		 dct[0][0] = cos00_term_quantized[31:0];
		 dct[0][1] = cos01_term_quantized[31:0];
		 dct[0][2] = cos02_term_quantized[31:0];
		 dct[0][3] = cos03_term_quantized[31:0];
		 dct[0][4] = cos04_term_quantized[31:0];
		 dct[0][5] = cos05_term_quantized[31:0];
		 dct[0][6] = cos06_term_quantized[31:0];
		 dct[0][7] = cos07_term_quantized[31:0];
		 dct[1][0] = cos10_term_quantized[31:0];
		 dct[1][1] = cos11_term_quantized[31:0];
		 dct[1][2] = cos12_term_quantized[31:0];
		 dct[1][3] = cos13_term_quantized[31:0];
		 dct[1][4] = cos14_term_quantized[31:0];
		 dct[1][5] = cos15_term_quantized[31:0];
		 dct[1][6] = cos16_term_quantized[31:0];
		 dct[1][7] = cos17_term_quantized[31:0];
		 dct[2][0] = cos20_term_quantized[31:0];
		 dct[2][1] = cos21_term_quantized[31:0];
		 dct[2][2] = cos22_term_quantized[31:0];
		 dct[2][3] = cos23_term_quantized[31:0];
		 dct[2][4] = cos24_term_quantized[31:0];
		 dct[2][5] = cos25_term_quantized[31:0];
		 dct[2][6] = cos26_term_quantized[31:0];
		 dct[2][7] = cos27_term_quantized[31:0];
		 dct[3][0] = cos30_term_quantized[31:0];
		 dct[3][1] = cos31_term_quantized[31:0];
		 dct[3][2] = cos32_term_quantized[31:0];
		 dct[3][3] = cos33_term_quantized[31:0];
		 dct[3][4] = cos34_term_quantized[31:0];
		 dct[3][5] = cos35_term_quantized[31:0];
		 dct[3][6] = cos36_term_quantized[31:0];
		 dct[3][7] = cos37_term_quantized[31:0];
		 dct[4][0] = cos40_term_quantized[31:0];
		 dct[4][1] = cos41_term_quantized[31:0];
		 dct[4][2] = cos42_term_quantized[31:0];
		 dct[4][3] = cos43_term_quantized[31:0];
		 dct[4][4] = cos44_term_quantized[31:0];
		 dct[4][5] = cos45_term_quantized[31:0];
		 dct[4][6] = cos46_term_quantized[31:0];
		 dct[4][7] = cos47_term_quantized[31:0];
		 dct[5][0] = cos50_term_quantized[31:0];
		 dct[5][1] = cos51_term_quantized[31:0];
		 dct[5][2] = cos52_term_quantized[31:0];
		 dct[5][3] = cos53_term_quantized[31:0];
		 dct[5][4] = cos54_term_quantized[31:0];
		 dct[5][5] = cos55_term_quantized[31:0];
		 dct[5][6] = cos56_term_quantized[31:0];
		 dct[5][7] = cos57_term_quantized[31:0];
		 dct[6][0] = cos60_term_quantized[31:0];
		 dct[6][1] = cos61_term_quantized[31:0];
		 dct[6][2] = cos62_term_quantized[31:0];
		 dct[6][3] = cos63_term_quantized[31:0];
		 dct[6][4] = cos64_term_quantized[31:0];
		 dct[6][5] = cos65_term_quantized[31:0];
		 dct[6][6] = cos66_term_quantized[31:0];
		 dct[6][7] = cos67_term_quantized[31:0];
		 dct[7][0] = cos70_term_quantized[31:0];
		 dct[7][1] = cos71_term_quantized[31:0];
		 dct[7][2] = cos72_term_quantized[31:0];
		 dct[7][3] = cos73_term_quantized[31:0];
		 dct[7][4] = cos74_term_quantized[31:0];
		 dct[7][5] = cos75_term_quantized[31:0];
		 dct[7][6] = cos76_term_quantized[31:0];
		 dct[7][7] = cos77_term_quantized[31:0];
	end
endmodule