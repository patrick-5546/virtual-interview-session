module dct_quantization(input logic [511:0] mcu, output logic [511:0] dct);
	wire[15:0] cos00_term = mcu[7:0] + mcu[15:8] + mcu[23:16] + mcu[31:24] + mcu[39:32] + mcu[47:40] + mcu[55:48] + mcu[63:56] + mcu[71:64] + mcu[79:72] + mcu[87:80] + mcu[95:88] + mcu[103:96] + mcu[111:104] + mcu[119:112] + mcu[127:120] + mcu[135:128] + mcu[143:136] + mcu[151:144] + mcu[159:152] + mcu[167:160] + mcu[175:168] + mcu[183:176] + mcu[191:184] + mcu[199:192] + mcu[207:200] + mcu[215:208] + mcu[223:216] + mcu[231:224] + mcu[239:232] + mcu[247:240] + mcu[255:248] + mcu[263:256] + mcu[271:264] + mcu[279:272] + mcu[287:280] + mcu[295:288] + mcu[303:296] + mcu[311:304] + mcu[319:312] + mcu[327:320] + mcu[335:328] + mcu[343:336] + mcu[351:344] + mcu[359:352] + mcu[367:360] + mcu[375:368] + mcu[383:376] + mcu[391:384] + mcu[399:392] + mcu[407:400] + mcu[415:408] + mcu[423:416] + mcu[431:424] + mcu[439:432] + mcu[447:440] + mcu[455:448] + mcu[463:456] + mcu[471:464] + mcu[479:472] + mcu[487:480] + mcu[495:488] + mcu[503:496] + mcu[511:504];
	wire[23:0] cos01_term = mcu[7:0] * 24'h0fb + mcu[15:8] * 24'h0d4 + mcu[23:16] * 24'h08e + mcu[31:24] * 24'h031 + mcu[39:32] * -24'h031 + mcu[47:40] * -24'h08e + mcu[55:48] * -24'h0d4 + mcu[63:56] * -24'h0fb + mcu[71:64] * 24'h0fb + mcu[79:72] * 24'h0d4 + mcu[87:80] * 24'h08e + mcu[95:88] * 24'h031 + mcu[103:96] * -24'h031 + mcu[111:104] * -24'h08e + mcu[119:112] * -24'h0d4 + mcu[127:120] * -24'h0fb + mcu[135:128] * 24'h0fb + mcu[143:136] * 24'h0d4 + mcu[151:144] * 24'h08e + mcu[159:152] * 24'h031 + mcu[167:160] * -24'h031 + mcu[175:168] * -24'h08e + mcu[183:176] * -24'h0d4 + mcu[191:184] * -24'h0fb + mcu[199:192] * 24'h0fb + mcu[207:200] * 24'h0d4 + mcu[215:208] * 24'h08e + mcu[223:216] * 24'h031 + mcu[231:224] * -24'h031 + mcu[239:232] * -24'h08e + mcu[247:240] * -24'h0d4 + mcu[255:248] * -24'h0fb + mcu[263:256] * 24'h0fb + mcu[271:264] * 24'h0d4 + mcu[279:272] * 24'h08e + mcu[287:280] * 24'h031 + mcu[295:288] * -24'h031 + mcu[303:296] * -24'h08e + mcu[311:304] * -24'h0d4 + mcu[319:312] * -24'h0fb + mcu[327:320] * 24'h0fb + mcu[335:328] * 24'h0d4 + mcu[343:336] * 24'h08e + mcu[351:344] * 24'h031 + mcu[359:352] * -24'h031 + mcu[367:360] * -24'h08e + mcu[375:368] * -24'h0d4 + mcu[383:376] * -24'h0fb + mcu[391:384] * 24'h0fb + mcu[399:392] * 24'h0d4 + mcu[407:400] * 24'h08e + mcu[415:408] * 24'h031 + mcu[423:416] * -24'h031 + mcu[431:424] * -24'h08e + mcu[439:432] * -24'h0d4 + mcu[447:440] * -24'h0fb + mcu[455:448] * 24'h0fb + mcu[463:456] * 24'h0d4 + mcu[471:464] * 24'h08e + mcu[479:472] * 24'h031 + mcu[487:480] * -24'h031 + mcu[495:488] * -24'h08e + mcu[503:496] * -24'h0d4 + mcu[511:504] * -24'h0fb;
	wire[23:0] cos02_term = mcu[7:0] * 24'h0ec + mcu[15:8] * 24'h062 + mcu[23:16] * -24'h062 + mcu[31:24] * -24'h0ec + mcu[39:32] * -24'h0ec + mcu[47:40] * -24'h062 + mcu[55:48] * 24'h062 + mcu[63:56] * 24'h0ec + mcu[71:64] * 24'h0ec + mcu[79:72] * 24'h062 + mcu[87:80] * -24'h062 + mcu[95:88] * -24'h0ec + mcu[103:96] * -24'h0ec + mcu[111:104] * -24'h062 + mcu[119:112] * 24'h062 + mcu[127:120] * 24'h0ec + mcu[135:128] * 24'h0ec + mcu[143:136] * 24'h062 + mcu[151:144] * -24'h062 + mcu[159:152] * -24'h0ec + mcu[167:160] * -24'h0ec + mcu[175:168] * -24'h062 + mcu[183:176] * 24'h062 + mcu[191:184] * 24'h0ec + mcu[199:192] * 24'h0ec + mcu[207:200] * 24'h062 + mcu[215:208] * -24'h062 + mcu[223:216] * -24'h0ec + mcu[231:224] * -24'h0ec + mcu[239:232] * -24'h062 + mcu[247:240] * 24'h062 + mcu[255:248] * 24'h0ec + mcu[263:256] * 24'h0ec + mcu[271:264] * 24'h062 + mcu[279:272] * -24'h062 + mcu[287:280] * -24'h0ec + mcu[295:288] * -24'h0ec + mcu[303:296] * -24'h062 + mcu[311:304] * 24'h062 + mcu[319:312] * 24'h0ec + mcu[327:320] * 24'h0ec + mcu[335:328] * 24'h062 + mcu[343:336] * -24'h062 + mcu[351:344] * -24'h0ec + mcu[359:352] * -24'h0ec + mcu[367:360] * -24'h062 + mcu[375:368] * 24'h062 + mcu[383:376] * 24'h0ec + mcu[391:384] * 24'h0ec + mcu[399:392] * 24'h062 + mcu[407:400] * -24'h062 + mcu[415:408] * -24'h0ec + mcu[423:416] * -24'h0ec + mcu[431:424] * -24'h062 + mcu[439:432] * 24'h062 + mcu[447:440] * 24'h0ec + mcu[455:448] * 24'h0ec + mcu[463:456] * 24'h062 + mcu[471:464] * -24'h062 + mcu[479:472] * -24'h0ec + mcu[487:480] * -24'h0ec + mcu[495:488] * -24'h062 + mcu[503:496] * 24'h062 + mcu[511:504] * 24'h0ec;
	wire[23:0] cos03_term = mcu[7:0] * 24'h0d4 + mcu[15:8] * -24'h031 + mcu[23:16] * -24'h0fb + mcu[31:24] * -24'h08e + mcu[39:32] * 24'h08e + mcu[47:40] * 24'h0fb + mcu[55:48] * 24'h031 + mcu[63:56] * -24'h0d4 + mcu[71:64] * 24'h0d4 + mcu[79:72] * -24'h031 + mcu[87:80] * -24'h0fb + mcu[95:88] * -24'h08e + mcu[103:96] * 24'h08e + mcu[111:104] * 24'h0fb + mcu[119:112] * 24'h031 + mcu[127:120] * -24'h0d4 + mcu[135:128] * 24'h0d4 + mcu[143:136] * -24'h031 + mcu[151:144] * -24'h0fb + mcu[159:152] * -24'h08e + mcu[167:160] * 24'h08e + mcu[175:168] * 24'h0fb + mcu[183:176] * 24'h031 + mcu[191:184] * -24'h0d4 + mcu[199:192] * 24'h0d4 + mcu[207:200] * -24'h031 + mcu[215:208] * -24'h0fb + mcu[223:216] * -24'h08e + mcu[231:224] * 24'h08e + mcu[239:232] * 24'h0fb + mcu[247:240] * 24'h031 + mcu[255:248] * -24'h0d4 + mcu[263:256] * 24'h0d4 + mcu[271:264] * -24'h031 + mcu[279:272] * -24'h0fb + mcu[287:280] * -24'h08e + mcu[295:288] * 24'h08e + mcu[303:296] * 24'h0fb + mcu[311:304] * 24'h031 + mcu[319:312] * -24'h0d4 + mcu[327:320] * 24'h0d4 + mcu[335:328] * -24'h031 + mcu[343:336] * -24'h0fb + mcu[351:344] * -24'h08e + mcu[359:352] * 24'h08e + mcu[367:360] * 24'h0fb + mcu[375:368] * 24'h031 + mcu[383:376] * -24'h0d4 + mcu[391:384] * 24'h0d4 + mcu[399:392] * -24'h031 + mcu[407:400] * -24'h0fb + mcu[415:408] * -24'h08e + mcu[423:416] * 24'h08e + mcu[431:424] * 24'h0fb + mcu[439:432] * 24'h031 + mcu[447:440] * -24'h0d4 + mcu[455:448] * 24'h0d4 + mcu[463:456] * -24'h031 + mcu[471:464] * -24'h0fb + mcu[479:472] * -24'h08e + mcu[487:480] * 24'h08e + mcu[495:488] * 24'h0fb + mcu[503:496] * 24'h031 + mcu[511:504] * -24'h0d4;
	wire[23:0] cos04_term = mcu[7:0] * 24'h0b4 + mcu[15:8] * -24'h0b4 + mcu[23:16] * -24'h0b4 + mcu[31:24] * 24'h0b4 + mcu[39:32] * 24'h0b4 + mcu[47:40] * -24'h0b4 + mcu[55:48] * -24'h0b4 + mcu[63:56] * 24'h0b4 + mcu[71:64] * 24'h0b4 + mcu[79:72] * -24'h0b4 + mcu[87:80] * -24'h0b4 + mcu[95:88] * 24'h0b4 + mcu[103:96] * 24'h0b4 + mcu[111:104] * -24'h0b4 + mcu[119:112] * -24'h0b4 + mcu[127:120] * 24'h0b4 + mcu[135:128] * 24'h0b4 + mcu[143:136] * -24'h0b4 + mcu[151:144] * -24'h0b4 + mcu[159:152] * 24'h0b4 + mcu[167:160] * 24'h0b4 + mcu[175:168] * -24'h0b4 + mcu[183:176] * -24'h0b4 + mcu[191:184] * 24'h0b4 + mcu[199:192] * 24'h0b4 + mcu[207:200] * -24'h0b4 + mcu[215:208] * -24'h0b4 + mcu[223:216] * 24'h0b4 + mcu[231:224] * 24'h0b4 + mcu[239:232] * -24'h0b4 + mcu[247:240] * -24'h0b4 + mcu[255:248] * 24'h0b4 + mcu[263:256] * 24'h0b4 + mcu[271:264] * -24'h0b4 + mcu[279:272] * -24'h0b4 + mcu[287:280] * 24'h0b4 + mcu[295:288] * 24'h0b4 + mcu[303:296] * -24'h0b4 + mcu[311:304] * -24'h0b4 + mcu[319:312] * 24'h0b4 + mcu[327:320] * 24'h0b4 + mcu[335:328] * -24'h0b4 + mcu[343:336] * -24'h0b4 + mcu[351:344] * 24'h0b4 + mcu[359:352] * 24'h0b4 + mcu[367:360] * -24'h0b4 + mcu[375:368] * -24'h0b4 + mcu[383:376] * 24'h0b4 + mcu[391:384] * 24'h0b4 + mcu[399:392] * -24'h0b4 + mcu[407:400] * -24'h0b4 + mcu[415:408] * 24'h0b4 + mcu[423:416] * 24'h0b4 + mcu[431:424] * -24'h0b4 + mcu[439:432] * -24'h0b4 + mcu[447:440] * 24'h0b4 + mcu[455:448] * 24'h0b4 + mcu[463:456] * -24'h0b4 + mcu[471:464] * -24'h0b4 + mcu[479:472] * 24'h0b4 + mcu[487:480] * 24'h0b4 + mcu[495:488] * -24'h0b4 + mcu[503:496] * -24'h0b4 + mcu[511:504] * 24'h0b4;
	wire[23:0] cos05_term = mcu[7:0] * 24'h08e + mcu[15:8] * -24'h0fb + mcu[23:16] * 24'h031 + mcu[31:24] * 24'h0d4 + mcu[39:32] * -24'h0d4 + mcu[47:40] * -24'h031 + mcu[55:48] * 24'h0fb + mcu[63:56] * -24'h08e + mcu[71:64] * 24'h08e + mcu[79:72] * -24'h0fb + mcu[87:80] * 24'h031 + mcu[95:88] * 24'h0d4 + mcu[103:96] * -24'h0d4 + mcu[111:104] * -24'h031 + mcu[119:112] * 24'h0fb + mcu[127:120] * -24'h08e + mcu[135:128] * 24'h08e + mcu[143:136] * -24'h0fb + mcu[151:144] * 24'h031 + mcu[159:152] * 24'h0d4 + mcu[167:160] * -24'h0d4 + mcu[175:168] * -24'h031 + mcu[183:176] * 24'h0fb + mcu[191:184] * -24'h08e + mcu[199:192] * 24'h08e + mcu[207:200] * -24'h0fb + mcu[215:208] * 24'h031 + mcu[223:216] * 24'h0d4 + mcu[231:224] * -24'h0d4 + mcu[239:232] * -24'h031 + mcu[247:240] * 24'h0fb + mcu[255:248] * -24'h08e + mcu[263:256] * 24'h08e + mcu[271:264] * -24'h0fb + mcu[279:272] * 24'h031 + mcu[287:280] * 24'h0d4 + mcu[295:288] * -24'h0d4 + mcu[303:296] * -24'h031 + mcu[311:304] * 24'h0fb + mcu[319:312] * -24'h08e + mcu[327:320] * 24'h08e + mcu[335:328] * -24'h0fb + mcu[343:336] * 24'h031 + mcu[351:344] * 24'h0d4 + mcu[359:352] * -24'h0d4 + mcu[367:360] * -24'h031 + mcu[375:368] * 24'h0fb + mcu[383:376] * -24'h08e + mcu[391:384] * 24'h08e + mcu[399:392] * -24'h0fb + mcu[407:400] * 24'h031 + mcu[415:408] * 24'h0d4 + mcu[423:416] * -24'h0d4 + mcu[431:424] * -24'h031 + mcu[439:432] * 24'h0fb + mcu[447:440] * -24'h08e + mcu[455:448] * 24'h08e + mcu[463:456] * -24'h0fb + mcu[471:464] * 24'h031 + mcu[479:472] * 24'h0d4 + mcu[487:480] * -24'h0d4 + mcu[495:488] * -24'h031 + mcu[503:496] * 24'h0fb + mcu[511:504] * -24'h08e;
	wire[23:0] cos06_term = mcu[7:0] * 24'h062 + mcu[15:8] * -24'h0ec + mcu[23:16] * 24'h0ec + mcu[31:24] * -24'h062 + mcu[39:32] * -24'h062 + mcu[47:40] * 24'h0ec + mcu[55:48] * -24'h0ec + mcu[63:56] * 24'h062 + mcu[71:64] * 24'h062 + mcu[79:72] * -24'h0ec + mcu[87:80] * 24'h0ec + mcu[95:88] * -24'h062 + mcu[103:96] * -24'h062 + mcu[111:104] * 24'h0ec + mcu[119:112] * -24'h0ec + mcu[127:120] * 24'h062 + mcu[135:128] * 24'h062 + mcu[143:136] * -24'h0ec + mcu[151:144] * 24'h0ec + mcu[159:152] * -24'h062 + mcu[167:160] * -24'h062 + mcu[175:168] * 24'h0ec + mcu[183:176] * -24'h0ec + mcu[191:184] * 24'h062 + mcu[199:192] * 24'h062 + mcu[207:200] * -24'h0ec + mcu[215:208] * 24'h0ec + mcu[223:216] * -24'h062 + mcu[231:224] * -24'h062 + mcu[239:232] * 24'h0ec + mcu[247:240] * -24'h0ec + mcu[255:248] * 24'h062 + mcu[263:256] * 24'h062 + mcu[271:264] * -24'h0ec + mcu[279:272] * 24'h0ec + mcu[287:280] * -24'h062 + mcu[295:288] * -24'h062 + mcu[303:296] * 24'h0ec + mcu[311:304] * -24'h0ec + mcu[319:312] * 24'h062 + mcu[327:320] * 24'h062 + mcu[335:328] * -24'h0ec + mcu[343:336] * 24'h0ec + mcu[351:344] * -24'h062 + mcu[359:352] * -24'h062 + mcu[367:360] * 24'h0ec + mcu[375:368] * -24'h0ec + mcu[383:376] * 24'h062 + mcu[391:384] * 24'h062 + mcu[399:392] * -24'h0ec + mcu[407:400] * 24'h0ec + mcu[415:408] * -24'h062 + mcu[423:416] * -24'h062 + mcu[431:424] * 24'h0ec + mcu[439:432] * -24'h0ec + mcu[447:440] * 24'h062 + mcu[455:448] * 24'h062 + mcu[463:456] * -24'h0ec + mcu[471:464] * 24'h0ec + mcu[479:472] * -24'h062 + mcu[487:480] * -24'h062 + mcu[495:488] * 24'h0ec + mcu[503:496] * -24'h0ec + mcu[511:504] * 24'h062;
	wire[23:0] cos07_term = mcu[7:0] * 24'h031 + mcu[15:8] * -24'h08e + mcu[23:16] * 24'h0d4 + mcu[31:24] * -24'h0fb + mcu[39:32] * 24'h0fb + mcu[47:40] * -24'h0d4 + mcu[55:48] * 24'h08e + mcu[63:56] * -24'h031 + mcu[71:64] * 24'h031 + mcu[79:72] * -24'h08e + mcu[87:80] * 24'h0d4 + mcu[95:88] * -24'h0fb + mcu[103:96] * 24'h0fb + mcu[111:104] * -24'h0d4 + mcu[119:112] * 24'h08e + mcu[127:120] * -24'h031 + mcu[135:128] * 24'h031 + mcu[143:136] * -24'h08e + mcu[151:144] * 24'h0d4 + mcu[159:152] * -24'h0fb + mcu[167:160] * 24'h0fb + mcu[175:168] * -24'h0d4 + mcu[183:176] * 24'h08e + mcu[191:184] * -24'h031 + mcu[199:192] * 24'h031 + mcu[207:200] * -24'h08e + mcu[215:208] * 24'h0d4 + mcu[223:216] * -24'h0fb + mcu[231:224] * 24'h0fb + mcu[239:232] * -24'h0d4 + mcu[247:240] * 24'h08e + mcu[255:248] * -24'h031 + mcu[263:256] * 24'h031 + mcu[271:264] * -24'h08e + mcu[279:272] * 24'h0d4 + mcu[287:280] * -24'h0fb + mcu[295:288] * 24'h0fb + mcu[303:296] * -24'h0d4 + mcu[311:304] * 24'h08e + mcu[319:312] * -24'h031 + mcu[327:320] * 24'h031 + mcu[335:328] * -24'h08e + mcu[343:336] * 24'h0d4 + mcu[351:344] * -24'h0fb + mcu[359:352] * 24'h0fb + mcu[367:360] * -24'h0d4 + mcu[375:368] * 24'h08e + mcu[383:376] * -24'h031 + mcu[391:384] * 24'h031 + mcu[399:392] * -24'h08e + mcu[407:400] * 24'h0d4 + mcu[415:408] * -24'h0fb + mcu[423:416] * 24'h0fb + mcu[431:424] * -24'h0d4 + mcu[439:432] * 24'h08e + mcu[447:440] * -24'h031 + mcu[455:448] * 24'h031 + mcu[463:456] * -24'h08e + mcu[471:464] * 24'h0d4 + mcu[479:472] * -24'h0fb + mcu[487:480] * 24'h0fb + mcu[495:488] * -24'h0d4 + mcu[503:496] * 24'h08e + mcu[511:504] * -24'h031;
	wire[23:0] cos10_term = mcu[7:0] * 24'h0fb + mcu[15:8] * 24'h0fb + mcu[23:16] * 24'h0fb + mcu[31:24] * 24'h0fb + mcu[39:32] * 24'h0fb + mcu[47:40] * 24'h0fb + mcu[55:48] * 24'h0fb + mcu[63:56] * 24'h0fb + mcu[71:64] * 24'h0d4 + mcu[79:72] * 24'h0d4 + mcu[87:80] * 24'h0d4 + mcu[95:88] * 24'h0d4 + mcu[103:96] * 24'h0d4 + mcu[111:104] * 24'h0d4 + mcu[119:112] * 24'h0d4 + mcu[127:120] * 24'h0d4 + mcu[135:128] * 24'h08e + mcu[143:136] * 24'h08e + mcu[151:144] * 24'h08e + mcu[159:152] * 24'h08e + mcu[167:160] * 24'h08e + mcu[175:168] * 24'h08e + mcu[183:176] * 24'h08e + mcu[191:184] * 24'h08e + mcu[199:192] * 24'h031 + mcu[207:200] * 24'h031 + mcu[215:208] * 24'h031 + mcu[223:216] * 24'h031 + mcu[231:224] * 24'h031 + mcu[239:232] * 24'h031 + mcu[247:240] * 24'h031 + mcu[255:248] * 24'h031 + mcu[263:256] * -24'h031 + mcu[271:264] * -24'h031 + mcu[279:272] * -24'h031 + mcu[287:280] * -24'h031 + mcu[295:288] * -24'h031 + mcu[303:296] * -24'h031 + mcu[311:304] * -24'h031 + mcu[319:312] * -24'h031 + mcu[327:320] * -24'h08e + mcu[335:328] * -24'h08e + mcu[343:336] * -24'h08e + mcu[351:344] * -24'h08e + mcu[359:352] * -24'h08e + mcu[367:360] * -24'h08e + mcu[375:368] * -24'h08e + mcu[383:376] * -24'h08e + mcu[391:384] * -24'h0d4 + mcu[399:392] * -24'h0d4 + mcu[407:400] * -24'h0d4 + mcu[415:408] * -24'h0d4 + mcu[423:416] * -24'h0d4 + mcu[431:424] * -24'h0d4 + mcu[439:432] * -24'h0d4 + mcu[447:440] * -24'h0d4 + mcu[455:448] * -24'h0fb + mcu[463:456] * -24'h0fb + mcu[471:464] * -24'h0fb + mcu[479:472] * -24'h0fb + mcu[487:480] * -24'h0fb + mcu[495:488] * -24'h0fb + mcu[503:496] * -24'h0fb + mcu[511:504] * -24'h0fb;
	wire[23:0] cos11_term = mcu[7:0] * 24'h0f6 + mcu[15:8] * 24'h0d0 + mcu[23:16] * 24'h08b + mcu[31:24] * 24'h030 + mcu[39:32] * -24'h030 + mcu[47:40] * -24'h08b + mcu[55:48] * -24'h0d0 + mcu[63:56] * -24'h0f6 + mcu[71:64] * 24'h0d0 + mcu[79:72] * 24'h0b0 + mcu[87:80] * 24'h076 + mcu[95:88] * 24'h029 + mcu[103:96] * -24'h029 + mcu[111:104] * -24'h076 + mcu[119:112] * -24'h0b0 + mcu[127:120] * -24'h0d0 + mcu[135:128] * 24'h08b + mcu[143:136] * 24'h076 + mcu[151:144] * 24'h04f + mcu[159:152] * 24'h01b + mcu[167:160] * -24'h01b + mcu[175:168] * -24'h04f + mcu[183:176] * -24'h076 + mcu[191:184] * -24'h08b + mcu[199:192] * 24'h030 + mcu[207:200] * 24'h029 + mcu[215:208] * 24'h01b + mcu[223:216] * 24'h009 + mcu[231:224] * -24'h009 + mcu[239:232] * -24'h01b + mcu[247:240] * -24'h029 + mcu[255:248] * -24'h030 + mcu[263:256] * -24'h030 + mcu[271:264] * -24'h029 + mcu[279:272] * -24'h01b + mcu[287:280] * -24'h009 + mcu[295:288] * 24'h009 + mcu[303:296] * 24'h01b + mcu[311:304] * 24'h029 + mcu[319:312] * 24'h030 + mcu[327:320] * -24'h08b + mcu[335:328] * -24'h076 + mcu[343:336] * -24'h04f + mcu[351:344] * -24'h01b + mcu[359:352] * 24'h01b + mcu[367:360] * 24'h04f + mcu[375:368] * 24'h076 + mcu[383:376] * 24'h08b + mcu[391:384] * -24'h0d0 + mcu[399:392] * -24'h0b0 + mcu[407:400] * -24'h076 + mcu[415:408] * -24'h029 + mcu[423:416] * 24'h029 + mcu[431:424] * 24'h076 + mcu[439:432] * 24'h0b0 + mcu[447:440] * 24'h0d0 + mcu[455:448] * -24'h0f6 + mcu[463:456] * -24'h0d0 + mcu[471:464] * -24'h08b + mcu[479:472] * -24'h030 + mcu[487:480] * 24'h030 + mcu[495:488] * 24'h08b + mcu[503:496] * 24'h0d0 + mcu[511:504] * 24'h0f6;
	wire[23:0] cos12_term = mcu[7:0] * 24'h0e7 + mcu[15:8] * 24'h060 + mcu[23:16] * -24'h060 + mcu[31:24] * -24'h0e7 + mcu[39:32] * -24'h0e7 + mcu[47:40] * -24'h060 + mcu[55:48] * 24'h060 + mcu[63:56] * 24'h0e7 + mcu[71:64] * 24'h0c4 + mcu[79:72] * 24'h051 + mcu[87:80] * -24'h051 + mcu[95:88] * -24'h0c4 + mcu[103:96] * -24'h0c4 + mcu[111:104] * -24'h051 + mcu[119:112] * 24'h051 + mcu[127:120] * 24'h0c4 + mcu[135:128] * 24'h083 + mcu[143:136] * 24'h036 + mcu[151:144] * -24'h036 + mcu[159:152] * -24'h083 + mcu[167:160] * -24'h083 + mcu[175:168] * -24'h036 + mcu[183:176] * 24'h036 + mcu[191:184] * 24'h083 + mcu[199:192] * 24'h02e + mcu[207:200] * 24'h013 + mcu[215:208] * -24'h013 + mcu[223:216] * -24'h02e + mcu[231:224] * -24'h02e + mcu[239:232] * -24'h013 + mcu[247:240] * 24'h013 + mcu[255:248] * 24'h02e + mcu[263:256] * -24'h02e + mcu[271:264] * -24'h013 + mcu[279:272] * 24'h013 + mcu[287:280] * 24'h02e + mcu[295:288] * 24'h02e + mcu[303:296] * 24'h013 + mcu[311:304] * -24'h013 + mcu[319:312] * -24'h02e + mcu[327:320] * -24'h083 + mcu[335:328] * -24'h036 + mcu[343:336] * 24'h036 + mcu[351:344] * 24'h083 + mcu[359:352] * 24'h083 + mcu[367:360] * 24'h036 + mcu[375:368] * -24'h036 + mcu[383:376] * -24'h083 + mcu[391:384] * -24'h0c4 + mcu[399:392] * -24'h051 + mcu[407:400] * 24'h051 + mcu[415:408] * 24'h0c4 + mcu[423:416] * 24'h0c4 + mcu[431:424] * 24'h051 + mcu[439:432] * -24'h051 + mcu[447:440] * -24'h0c4 + mcu[455:448] * -24'h0e7 + mcu[463:456] * -24'h060 + mcu[471:464] * 24'h060 + mcu[479:472] * 24'h0e7 + mcu[487:480] * 24'h0e7 + mcu[495:488] * 24'h060 + mcu[503:496] * -24'h060 + mcu[511:504] * -24'h0e7;
	wire[23:0] cos13_term = mcu[7:0] * 24'h0d0 + mcu[15:8] * -24'h030 + mcu[23:16] * -24'h0f6 + mcu[31:24] * -24'h08b + mcu[39:32] * 24'h08b + mcu[47:40] * 24'h0f6 + mcu[55:48] * 24'h030 + mcu[63:56] * -24'h0d0 + mcu[71:64] * 24'h0b0 + mcu[79:72] * -24'h029 + mcu[87:80] * -24'h0d0 + mcu[95:88] * -24'h076 + mcu[103:96] * 24'h076 + mcu[111:104] * 24'h0d0 + mcu[119:112] * 24'h029 + mcu[127:120] * -24'h0b0 + mcu[135:128] * 24'h076 + mcu[143:136] * -24'h01b + mcu[151:144] * -24'h08b + mcu[159:152] * -24'h04f + mcu[167:160] * 24'h04f + mcu[175:168] * 24'h08b + mcu[183:176] * 24'h01b + mcu[191:184] * -24'h076 + mcu[199:192] * 24'h029 + mcu[207:200] * -24'h009 + mcu[215:208] * -24'h030 + mcu[223:216] * -24'h01b + mcu[231:224] * 24'h01b + mcu[239:232] * 24'h030 + mcu[247:240] * 24'h009 + mcu[255:248] * -24'h029 + mcu[263:256] * -24'h029 + mcu[271:264] * 24'h009 + mcu[279:272] * 24'h030 + mcu[287:280] * 24'h01b + mcu[295:288] * -24'h01b + mcu[303:296] * -24'h030 + mcu[311:304] * -24'h009 + mcu[319:312] * 24'h029 + mcu[327:320] * -24'h076 + mcu[335:328] * 24'h01b + mcu[343:336] * 24'h08b + mcu[351:344] * 24'h04f + mcu[359:352] * -24'h04f + mcu[367:360] * -24'h08b + mcu[375:368] * -24'h01b + mcu[383:376] * 24'h076 + mcu[391:384] * -24'h0b0 + mcu[399:392] * 24'h029 + mcu[407:400] * 24'h0d0 + mcu[415:408] * 24'h076 + mcu[423:416] * -24'h076 + mcu[431:424] * -24'h0d0 + mcu[439:432] * -24'h029 + mcu[447:440] * 24'h0b0 + mcu[455:448] * -24'h0d0 + mcu[463:456] * 24'h030 + mcu[471:464] * 24'h0f6 + mcu[479:472] * 24'h08b + mcu[487:480] * -24'h08b + mcu[495:488] * -24'h0f6 + mcu[503:496] * -24'h030 + mcu[511:504] * 24'h0d0;
	wire[23:0] cos14_term = mcu[7:0] * 24'h0b1 + mcu[15:8] * -24'h0b1 + mcu[23:16] * -24'h0b1 + mcu[31:24] * 24'h0b1 + mcu[39:32] * 24'h0b1 + mcu[47:40] * -24'h0b1 + mcu[55:48] * -24'h0b1 + mcu[63:56] * 24'h0b1 + mcu[71:64] * 24'h096 + mcu[79:72] * -24'h096 + mcu[87:80] * -24'h096 + mcu[95:88] * 24'h096 + mcu[103:96] * 24'h096 + mcu[111:104] * -24'h096 + mcu[119:112] * -24'h096 + mcu[127:120] * 24'h096 + mcu[135:128] * 24'h064 + mcu[143:136] * -24'h064 + mcu[151:144] * -24'h064 + mcu[159:152] * 24'h064 + mcu[167:160] * 24'h064 + mcu[175:168] * -24'h064 + mcu[183:176] * -24'h064 + mcu[191:184] * 24'h064 + mcu[199:192] * 24'h023 + mcu[207:200] * -24'h023 + mcu[215:208] * -24'h023 + mcu[223:216] * 24'h023 + mcu[231:224] * 24'h023 + mcu[239:232] * -24'h023 + mcu[247:240] * -24'h023 + mcu[255:248] * 24'h023 + mcu[263:256] * -24'h023 + mcu[271:264] * 24'h023 + mcu[279:272] * 24'h023 + mcu[287:280] * -24'h023 + mcu[295:288] * -24'h023 + mcu[303:296] * 24'h023 + mcu[311:304] * 24'h023 + mcu[319:312] * -24'h023 + mcu[327:320] * -24'h064 + mcu[335:328] * 24'h064 + mcu[343:336] * 24'h064 + mcu[351:344] * -24'h064 + mcu[359:352] * -24'h064 + mcu[367:360] * 24'h064 + mcu[375:368] * 24'h064 + mcu[383:376] * -24'h064 + mcu[391:384] * -24'h096 + mcu[399:392] * 24'h096 + mcu[407:400] * 24'h096 + mcu[415:408] * -24'h096 + mcu[423:416] * -24'h096 + mcu[431:424] * 24'h096 + mcu[439:432] * 24'h096 + mcu[447:440] * -24'h096 + mcu[455:448] * -24'h0b1 + mcu[463:456] * 24'h0b1 + mcu[471:464] * 24'h0b1 + mcu[479:472] * -24'h0b1 + mcu[487:480] * -24'h0b1 + mcu[495:488] * 24'h0b1 + mcu[503:496] * 24'h0b1 + mcu[511:504] * -24'h0b1;
	wire[23:0] cos15_term = mcu[7:0] * 24'h08b + mcu[15:8] * -24'h0f6 + mcu[23:16] * 24'h030 + mcu[31:24] * 24'h0d0 + mcu[39:32] * -24'h0d0 + mcu[47:40] * -24'h030 + mcu[55:48] * 24'h0f6 + mcu[63:56] * -24'h08b + mcu[71:64] * 24'h076 + mcu[79:72] * -24'h0d0 + mcu[87:80] * 24'h029 + mcu[95:88] * 24'h0b0 + mcu[103:96] * -24'h0b0 + mcu[111:104] * -24'h029 + mcu[119:112] * 24'h0d0 + mcu[127:120] * -24'h076 + mcu[135:128] * 24'h04f + mcu[143:136] * -24'h08b + mcu[151:144] * 24'h01b + mcu[159:152] * 24'h076 + mcu[167:160] * -24'h076 + mcu[175:168] * -24'h01b + mcu[183:176] * 24'h08b + mcu[191:184] * -24'h04f + mcu[199:192] * 24'h01b + mcu[207:200] * -24'h030 + mcu[215:208] * 24'h009 + mcu[223:216] * 24'h029 + mcu[231:224] * -24'h029 + mcu[239:232] * -24'h009 + mcu[247:240] * 24'h030 + mcu[255:248] * -24'h01b + mcu[263:256] * -24'h01b + mcu[271:264] * 24'h030 + mcu[279:272] * -24'h009 + mcu[287:280] * -24'h029 + mcu[295:288] * 24'h029 + mcu[303:296] * 24'h009 + mcu[311:304] * -24'h030 + mcu[319:312] * 24'h01b + mcu[327:320] * -24'h04f + mcu[335:328] * 24'h08b + mcu[343:336] * -24'h01b + mcu[351:344] * -24'h076 + mcu[359:352] * 24'h076 + mcu[367:360] * 24'h01b + mcu[375:368] * -24'h08b + mcu[383:376] * 24'h04f + mcu[391:384] * -24'h076 + mcu[399:392] * 24'h0d0 + mcu[407:400] * -24'h029 + mcu[415:408] * -24'h0b0 + mcu[423:416] * 24'h0b0 + mcu[431:424] * 24'h029 + mcu[439:432] * -24'h0d0 + mcu[447:440] * 24'h076 + mcu[455:448] * -24'h08b + mcu[463:456] * 24'h0f6 + mcu[471:464] * -24'h030 + mcu[479:472] * -24'h0d0 + mcu[487:480] * 24'h0d0 + mcu[495:488] * 24'h030 + mcu[503:496] * -24'h0f6 + mcu[511:504] * 24'h08b;
	wire[23:0] cos16_term = mcu[7:0] * 24'h060 + mcu[15:8] * -24'h0e7 + mcu[23:16] * 24'h0e7 + mcu[31:24] * -24'h060 + mcu[39:32] * -24'h060 + mcu[47:40] * 24'h0e7 + mcu[55:48] * -24'h0e7 + mcu[63:56] * 24'h060 + mcu[71:64] * 24'h051 + mcu[79:72] * -24'h0c4 + mcu[87:80] * 24'h0c4 + mcu[95:88] * -24'h051 + mcu[103:96] * -24'h051 + mcu[111:104] * 24'h0c4 + mcu[119:112] * -24'h0c4 + mcu[127:120] * 24'h051 + mcu[135:128] * 24'h036 + mcu[143:136] * -24'h083 + mcu[151:144] * 24'h083 + mcu[159:152] * -24'h036 + mcu[167:160] * -24'h036 + mcu[175:168] * 24'h083 + mcu[183:176] * -24'h083 + mcu[191:184] * 24'h036 + mcu[199:192] * 24'h013 + mcu[207:200] * -24'h02e + mcu[215:208] * 24'h02e + mcu[223:216] * -24'h013 + mcu[231:224] * -24'h013 + mcu[239:232] * 24'h02e + mcu[247:240] * -24'h02e + mcu[255:248] * 24'h013 + mcu[263:256] * -24'h013 + mcu[271:264] * 24'h02e + mcu[279:272] * -24'h02e + mcu[287:280] * 24'h013 + mcu[295:288] * 24'h013 + mcu[303:296] * -24'h02e + mcu[311:304] * 24'h02e + mcu[319:312] * -24'h013 + mcu[327:320] * -24'h036 + mcu[335:328] * 24'h083 + mcu[343:336] * -24'h083 + mcu[351:344] * 24'h036 + mcu[359:352] * 24'h036 + mcu[367:360] * -24'h083 + mcu[375:368] * 24'h083 + mcu[383:376] * -24'h036 + mcu[391:384] * -24'h051 + mcu[399:392] * 24'h0c4 + mcu[407:400] * -24'h0c4 + mcu[415:408] * 24'h051 + mcu[423:416] * 24'h051 + mcu[431:424] * -24'h0c4 + mcu[439:432] * 24'h0c4 + mcu[447:440] * -24'h051 + mcu[455:448] * -24'h060 + mcu[463:456] * 24'h0e7 + mcu[471:464] * -24'h0e7 + mcu[479:472] * 24'h060 + mcu[487:480] * 24'h060 + mcu[495:488] * -24'h0e7 + mcu[503:496] * 24'h0e7 + mcu[511:504] * -24'h060;
	wire[23:0] cos17_term = mcu[7:0] * 24'h030 + mcu[15:8] * -24'h08b + mcu[23:16] * 24'h0d0 + mcu[31:24] * -24'h0f6 + mcu[39:32] * 24'h0f6 + mcu[47:40] * -24'h0d0 + mcu[55:48] * 24'h08b + mcu[63:56] * -24'h030 + mcu[71:64] * 24'h029 + mcu[79:72] * -24'h076 + mcu[87:80] * 24'h0b0 + mcu[95:88] * -24'h0d0 + mcu[103:96] * 24'h0d0 + mcu[111:104] * -24'h0b0 + mcu[119:112] * 24'h076 + mcu[127:120] * -24'h029 + mcu[135:128] * 24'h01b + mcu[143:136] * -24'h04f + mcu[151:144] * 24'h076 + mcu[159:152] * -24'h08b + mcu[167:160] * 24'h08b + mcu[175:168] * -24'h076 + mcu[183:176] * 24'h04f + mcu[191:184] * -24'h01b + mcu[199:192] * 24'h009 + mcu[207:200] * -24'h01b + mcu[215:208] * 24'h029 + mcu[223:216] * -24'h030 + mcu[231:224] * 24'h030 + mcu[239:232] * -24'h029 + mcu[247:240] * 24'h01b + mcu[255:248] * -24'h009 + mcu[263:256] * -24'h009 + mcu[271:264] * 24'h01b + mcu[279:272] * -24'h029 + mcu[287:280] * 24'h030 + mcu[295:288] * -24'h030 + mcu[303:296] * 24'h029 + mcu[311:304] * -24'h01b + mcu[319:312] * 24'h009 + mcu[327:320] * -24'h01b + mcu[335:328] * 24'h04f + mcu[343:336] * -24'h076 + mcu[351:344] * 24'h08b + mcu[359:352] * -24'h08b + mcu[367:360] * 24'h076 + mcu[375:368] * -24'h04f + mcu[383:376] * 24'h01b + mcu[391:384] * -24'h029 + mcu[399:392] * 24'h076 + mcu[407:400] * -24'h0b0 + mcu[415:408] * 24'h0d0 + mcu[423:416] * -24'h0d0 + mcu[431:424] * 24'h0b0 + mcu[439:432] * -24'h076 + mcu[447:440] * 24'h029 + mcu[455:448] * -24'h030 + mcu[463:456] * 24'h08b + mcu[471:464] * -24'h0d0 + mcu[479:472] * 24'h0f6 + mcu[487:480] * -24'h0f6 + mcu[495:488] * 24'h0d0 + mcu[503:496] * -24'h08b + mcu[511:504] * 24'h030;
	wire[23:0] cos20_term = mcu[7:0] * 24'h0ec + mcu[15:8] * 24'h0ec + mcu[23:16] * 24'h0ec + mcu[31:24] * 24'h0ec + mcu[39:32] * 24'h0ec + mcu[47:40] * 24'h0ec + mcu[55:48] * 24'h0ec + mcu[63:56] * 24'h0ec + mcu[71:64] * 24'h062 + mcu[79:72] * 24'h062 + mcu[87:80] * 24'h062 + mcu[95:88] * 24'h062 + mcu[103:96] * 24'h062 + mcu[111:104] * 24'h062 + mcu[119:112] * 24'h062 + mcu[127:120] * 24'h062 + mcu[135:128] * -24'h062 + mcu[143:136] * -24'h062 + mcu[151:144] * -24'h062 + mcu[159:152] * -24'h062 + mcu[167:160] * -24'h062 + mcu[175:168] * -24'h062 + mcu[183:176] * -24'h062 + mcu[191:184] * -24'h062 + mcu[199:192] * -24'h0ec + mcu[207:200] * -24'h0ec + mcu[215:208] * -24'h0ec + mcu[223:216] * -24'h0ec + mcu[231:224] * -24'h0ec + mcu[239:232] * -24'h0ec + mcu[247:240] * -24'h0ec + mcu[255:248] * -24'h0ec + mcu[263:256] * -24'h0ec + mcu[271:264] * -24'h0ec + mcu[279:272] * -24'h0ec + mcu[287:280] * -24'h0ec + mcu[295:288] * -24'h0ec + mcu[303:296] * -24'h0ec + mcu[311:304] * -24'h0ec + mcu[319:312] * -24'h0ec + mcu[327:320] * -24'h062 + mcu[335:328] * -24'h062 + mcu[343:336] * -24'h062 + mcu[351:344] * -24'h062 + mcu[359:352] * -24'h062 + mcu[367:360] * -24'h062 + mcu[375:368] * -24'h062 + mcu[383:376] * -24'h062 + mcu[391:384] * 24'h062 + mcu[399:392] * 24'h062 + mcu[407:400] * 24'h062 + mcu[415:408] * 24'h062 + mcu[423:416] * 24'h062 + mcu[431:424] * 24'h062 + mcu[439:432] * 24'h062 + mcu[447:440] * 24'h062 + mcu[455:448] * 24'h0ec + mcu[463:456] * 24'h0ec + mcu[471:464] * 24'h0ec + mcu[479:472] * 24'h0ec + mcu[487:480] * 24'h0ec + mcu[495:488] * 24'h0ec + mcu[503:496] * 24'h0ec + mcu[511:504] * 24'h0ec;
	wire[23:0] cos21_term = mcu[7:0] * 24'h0e7 + mcu[15:8] * 24'h0c4 + mcu[23:16] * 24'h083 + mcu[31:24] * 24'h02e + mcu[39:32] * -24'h02e + mcu[47:40] * -24'h083 + mcu[55:48] * -24'h0c4 + mcu[63:56] * -24'h0e7 + mcu[71:64] * 24'h060 + mcu[79:72] * 24'h051 + mcu[87:80] * 24'h036 + mcu[95:88] * 24'h013 + mcu[103:96] * -24'h013 + mcu[111:104] * -24'h036 + mcu[119:112] * -24'h051 + mcu[127:120] * -24'h060 + mcu[135:128] * -24'h060 + mcu[143:136] * -24'h051 + mcu[151:144] * -24'h036 + mcu[159:152] * -24'h013 + mcu[167:160] * 24'h013 + mcu[175:168] * 24'h036 + mcu[183:176] * 24'h051 + mcu[191:184] * 24'h060 + mcu[199:192] * -24'h0e7 + mcu[207:200] * -24'h0c4 + mcu[215:208] * -24'h083 + mcu[223:216] * -24'h02e + mcu[231:224] * 24'h02e + mcu[239:232] * 24'h083 + mcu[247:240] * 24'h0c4 + mcu[255:248] * 24'h0e7 + mcu[263:256] * -24'h0e7 + mcu[271:264] * -24'h0c4 + mcu[279:272] * -24'h083 + mcu[287:280] * -24'h02e + mcu[295:288] * 24'h02e + mcu[303:296] * 24'h083 + mcu[311:304] * 24'h0c4 + mcu[319:312] * 24'h0e7 + mcu[327:320] * -24'h060 + mcu[335:328] * -24'h051 + mcu[343:336] * -24'h036 + mcu[351:344] * -24'h013 + mcu[359:352] * 24'h013 + mcu[367:360] * 24'h036 + mcu[375:368] * 24'h051 + mcu[383:376] * 24'h060 + mcu[391:384] * 24'h060 + mcu[399:392] * 24'h051 + mcu[407:400] * 24'h036 + mcu[415:408] * 24'h013 + mcu[423:416] * -24'h013 + mcu[431:424] * -24'h036 + mcu[439:432] * -24'h051 + mcu[447:440] * -24'h060 + mcu[455:448] * 24'h0e7 + mcu[463:456] * 24'h0c4 + mcu[471:464] * 24'h083 + mcu[479:472] * 24'h02e + mcu[487:480] * -24'h02e + mcu[495:488] * -24'h083 + mcu[503:496] * -24'h0c4 + mcu[511:504] * -24'h0e7;
	wire[23:0] cos22_term = mcu[7:0] * 24'h0da + mcu[15:8] * 24'h05a + mcu[23:16] * -24'h05a + mcu[31:24] * -24'h0da + mcu[39:32] * -24'h0da + mcu[47:40] * -24'h05a + mcu[55:48] * 24'h05a + mcu[63:56] * 24'h0da + mcu[71:64] * 24'h05a + mcu[79:72] * 24'h025 + mcu[87:80] * -24'h025 + mcu[95:88] * -24'h05a + mcu[103:96] * -24'h05a + mcu[111:104] * -24'h025 + mcu[119:112] * 24'h025 + mcu[127:120] * 24'h05a + mcu[135:128] * -24'h05a + mcu[143:136] * -24'h025 + mcu[151:144] * 24'h025 + mcu[159:152] * 24'h05a + mcu[167:160] * 24'h05a + mcu[175:168] * 24'h025 + mcu[183:176] * -24'h025 + mcu[191:184] * -24'h05a + mcu[199:192] * -24'h0da + mcu[207:200] * -24'h05a + mcu[215:208] * 24'h05a + mcu[223:216] * 24'h0da + mcu[231:224] * 24'h0da + mcu[239:232] * 24'h05a + mcu[247:240] * -24'h05a + mcu[255:248] * -24'h0da + mcu[263:256] * -24'h0da + mcu[271:264] * -24'h05a + mcu[279:272] * 24'h05a + mcu[287:280] * 24'h0da + mcu[295:288] * 24'h0da + mcu[303:296] * 24'h05a + mcu[311:304] * -24'h05a + mcu[319:312] * -24'h0da + mcu[327:320] * -24'h05a + mcu[335:328] * -24'h025 + mcu[343:336] * 24'h025 + mcu[351:344] * 24'h05a + mcu[359:352] * 24'h05a + mcu[367:360] * 24'h025 + mcu[375:368] * -24'h025 + mcu[383:376] * -24'h05a + mcu[391:384] * 24'h05a + mcu[399:392] * 24'h025 + mcu[407:400] * -24'h025 + mcu[415:408] * -24'h05a + mcu[423:416] * -24'h05a + mcu[431:424] * -24'h025 + mcu[439:432] * 24'h025 + mcu[447:440] * 24'h05a + mcu[455:448] * 24'h0da + mcu[463:456] * 24'h05a + mcu[471:464] * -24'h05a + mcu[479:472] * -24'h0da + mcu[487:480] * -24'h0da + mcu[495:488] * -24'h05a + mcu[503:496] * 24'h05a + mcu[511:504] * 24'h0da;
	wire[23:0] cos23_term = mcu[7:0] * 24'h0c4 + mcu[15:8] * -24'h02e + mcu[23:16] * -24'h0e7 + mcu[31:24] * -24'h083 + mcu[39:32] * 24'h083 + mcu[47:40] * 24'h0e7 + mcu[55:48] * 24'h02e + mcu[63:56] * -24'h0c4 + mcu[71:64] * 24'h051 + mcu[79:72] * -24'h013 + mcu[87:80] * -24'h060 + mcu[95:88] * -24'h036 + mcu[103:96] * 24'h036 + mcu[111:104] * 24'h060 + mcu[119:112] * 24'h013 + mcu[127:120] * -24'h051 + mcu[135:128] * -24'h051 + mcu[143:136] * 24'h013 + mcu[151:144] * 24'h060 + mcu[159:152] * 24'h036 + mcu[167:160] * -24'h036 + mcu[175:168] * -24'h060 + mcu[183:176] * -24'h013 + mcu[191:184] * 24'h051 + mcu[199:192] * -24'h0c4 + mcu[207:200] * 24'h02e + mcu[215:208] * 24'h0e7 + mcu[223:216] * 24'h083 + mcu[231:224] * -24'h083 + mcu[239:232] * -24'h0e7 + mcu[247:240] * -24'h02e + mcu[255:248] * 24'h0c4 + mcu[263:256] * -24'h0c4 + mcu[271:264] * 24'h02e + mcu[279:272] * 24'h0e7 + mcu[287:280] * 24'h083 + mcu[295:288] * -24'h083 + mcu[303:296] * -24'h0e7 + mcu[311:304] * -24'h02e + mcu[319:312] * 24'h0c4 + mcu[327:320] * -24'h051 + mcu[335:328] * 24'h013 + mcu[343:336] * 24'h060 + mcu[351:344] * 24'h036 + mcu[359:352] * -24'h036 + mcu[367:360] * -24'h060 + mcu[375:368] * -24'h013 + mcu[383:376] * 24'h051 + mcu[391:384] * 24'h051 + mcu[399:392] * -24'h013 + mcu[407:400] * -24'h060 + mcu[415:408] * -24'h036 + mcu[423:416] * 24'h036 + mcu[431:424] * 24'h060 + mcu[439:432] * 24'h013 + mcu[447:440] * -24'h051 + mcu[455:448] * 24'h0c4 + mcu[463:456] * -24'h02e + mcu[471:464] * -24'h0e7 + mcu[479:472] * -24'h083 + mcu[487:480] * 24'h083 + mcu[495:488] * 24'h0e7 + mcu[503:496] * 24'h02e + mcu[511:504] * -24'h0c4;
	wire[23:0] cos24_term = mcu[7:0] * 24'h0a7 + mcu[15:8] * -24'h0a7 + mcu[23:16] * -24'h0a7 + mcu[31:24] * 24'h0a7 + mcu[39:32] * 24'h0a7 + mcu[47:40] * -24'h0a7 + mcu[55:48] * -24'h0a7 + mcu[63:56] * 24'h0a7 + mcu[71:64] * 24'h045 + mcu[79:72] * -24'h045 + mcu[87:80] * -24'h045 + mcu[95:88] * 24'h045 + mcu[103:96] * 24'h045 + mcu[111:104] * -24'h045 + mcu[119:112] * -24'h045 + mcu[127:120] * 24'h045 + mcu[135:128] * -24'h045 + mcu[143:136] * 24'h045 + mcu[151:144] * 24'h045 + mcu[159:152] * -24'h045 + mcu[167:160] * -24'h045 + mcu[175:168] * 24'h045 + mcu[183:176] * 24'h045 + mcu[191:184] * -24'h045 + mcu[199:192] * -24'h0a7 + mcu[207:200] * 24'h0a7 + mcu[215:208] * 24'h0a7 + mcu[223:216] * -24'h0a7 + mcu[231:224] * -24'h0a7 + mcu[239:232] * 24'h0a7 + mcu[247:240] * 24'h0a7 + mcu[255:248] * -24'h0a7 + mcu[263:256] * -24'h0a7 + mcu[271:264] * 24'h0a7 + mcu[279:272] * 24'h0a7 + mcu[287:280] * -24'h0a7 + mcu[295:288] * -24'h0a7 + mcu[303:296] * 24'h0a7 + mcu[311:304] * 24'h0a7 + mcu[319:312] * -24'h0a7 + mcu[327:320] * -24'h045 + mcu[335:328] * 24'h045 + mcu[343:336] * 24'h045 + mcu[351:344] * -24'h045 + mcu[359:352] * -24'h045 + mcu[367:360] * 24'h045 + mcu[375:368] * 24'h045 + mcu[383:376] * -24'h045 + mcu[391:384] * 24'h045 + mcu[399:392] * -24'h045 + mcu[407:400] * -24'h045 + mcu[415:408] * 24'h045 + mcu[423:416] * 24'h045 + mcu[431:424] * -24'h045 + mcu[439:432] * -24'h045 + mcu[447:440] * 24'h045 + mcu[455:448] * 24'h0a7 + mcu[463:456] * -24'h0a7 + mcu[471:464] * -24'h0a7 + mcu[479:472] * 24'h0a7 + mcu[487:480] * 24'h0a7 + mcu[495:488] * -24'h0a7 + mcu[503:496] * -24'h0a7 + mcu[511:504] * 24'h0a7;
	wire[23:0] cos25_term = mcu[7:0] * 24'h083 + mcu[15:8] * -24'h0e7 + mcu[23:16] * 24'h02e + mcu[31:24] * 24'h0c4 + mcu[39:32] * -24'h0c4 + mcu[47:40] * -24'h02e + mcu[55:48] * 24'h0e7 + mcu[63:56] * -24'h083 + mcu[71:64] * 24'h036 + mcu[79:72] * -24'h060 + mcu[87:80] * 24'h013 + mcu[95:88] * 24'h051 + mcu[103:96] * -24'h051 + mcu[111:104] * -24'h013 + mcu[119:112] * 24'h060 + mcu[127:120] * -24'h036 + mcu[135:128] * -24'h036 + mcu[143:136] * 24'h060 + mcu[151:144] * -24'h013 + mcu[159:152] * -24'h051 + mcu[167:160] * 24'h051 + mcu[175:168] * 24'h013 + mcu[183:176] * -24'h060 + mcu[191:184] * 24'h036 + mcu[199:192] * -24'h083 + mcu[207:200] * 24'h0e7 + mcu[215:208] * -24'h02e + mcu[223:216] * -24'h0c4 + mcu[231:224] * 24'h0c4 + mcu[239:232] * 24'h02e + mcu[247:240] * -24'h0e7 + mcu[255:248] * 24'h083 + mcu[263:256] * -24'h083 + mcu[271:264] * 24'h0e7 + mcu[279:272] * -24'h02e + mcu[287:280] * -24'h0c4 + mcu[295:288] * 24'h0c4 + mcu[303:296] * 24'h02e + mcu[311:304] * -24'h0e7 + mcu[319:312] * 24'h083 + mcu[327:320] * -24'h036 + mcu[335:328] * 24'h060 + mcu[343:336] * -24'h013 + mcu[351:344] * -24'h051 + mcu[359:352] * 24'h051 + mcu[367:360] * 24'h013 + mcu[375:368] * -24'h060 + mcu[383:376] * 24'h036 + mcu[391:384] * 24'h036 + mcu[399:392] * -24'h060 + mcu[407:400] * 24'h013 + mcu[415:408] * 24'h051 + mcu[423:416] * -24'h051 + mcu[431:424] * -24'h013 + mcu[439:432] * 24'h060 + mcu[447:440] * -24'h036 + mcu[455:448] * 24'h083 + mcu[463:456] * -24'h0e7 + mcu[471:464] * 24'h02e + mcu[479:472] * 24'h0c4 + mcu[487:480] * -24'h0c4 + mcu[495:488] * -24'h02e + mcu[503:496] * 24'h0e7 + mcu[511:504] * -24'h083;
	wire[23:0] cos26_term = mcu[7:0] * 24'h05a + mcu[15:8] * -24'h0da + mcu[23:16] * 24'h0da + mcu[31:24] * -24'h05a + mcu[39:32] * -24'h05a + mcu[47:40] * 24'h0da + mcu[55:48] * -24'h0da + mcu[63:56] * 24'h05a + mcu[71:64] * 24'h025 + mcu[79:72] * -24'h05a + mcu[87:80] * 24'h05a + mcu[95:88] * -24'h025 + mcu[103:96] * -24'h025 + mcu[111:104] * 24'h05a + mcu[119:112] * -24'h05a + mcu[127:120] * 24'h025 + mcu[135:128] * -24'h025 + mcu[143:136] * 24'h05a + mcu[151:144] * -24'h05a + mcu[159:152] * 24'h025 + mcu[167:160] * 24'h025 + mcu[175:168] * -24'h05a + mcu[183:176] * 24'h05a + mcu[191:184] * -24'h025 + mcu[199:192] * -24'h05a + mcu[207:200] * 24'h0da + mcu[215:208] * -24'h0da + mcu[223:216] * 24'h05a + mcu[231:224] * 24'h05a + mcu[239:232] * -24'h0da + mcu[247:240] * 24'h0da + mcu[255:248] * -24'h05a + mcu[263:256] * -24'h05a + mcu[271:264] * 24'h0da + mcu[279:272] * -24'h0da + mcu[287:280] * 24'h05a + mcu[295:288] * 24'h05a + mcu[303:296] * -24'h0da + mcu[311:304] * 24'h0da + mcu[319:312] * -24'h05a + mcu[327:320] * -24'h025 + mcu[335:328] * 24'h05a + mcu[343:336] * -24'h05a + mcu[351:344] * 24'h025 + mcu[359:352] * 24'h025 + mcu[367:360] * -24'h05a + mcu[375:368] * 24'h05a + mcu[383:376] * -24'h025 + mcu[391:384] * 24'h025 + mcu[399:392] * -24'h05a + mcu[407:400] * 24'h05a + mcu[415:408] * -24'h025 + mcu[423:416] * -24'h025 + mcu[431:424] * 24'h05a + mcu[439:432] * -24'h05a + mcu[447:440] * 24'h025 + mcu[455:448] * 24'h05a + mcu[463:456] * -24'h0da + mcu[471:464] * 24'h0da + mcu[479:472] * -24'h05a + mcu[487:480] * -24'h05a + mcu[495:488] * 24'h0da + mcu[503:496] * -24'h0da + mcu[511:504] * 24'h05a;
	wire[23:0] cos27_term = mcu[7:0] * 24'h02e + mcu[15:8] * -24'h083 + mcu[23:16] * 24'h0c4 + mcu[31:24] * -24'h0e7 + mcu[39:32] * 24'h0e7 + mcu[47:40] * -24'h0c4 + mcu[55:48] * 24'h083 + mcu[63:56] * -24'h02e + mcu[71:64] * 24'h013 + mcu[79:72] * -24'h036 + mcu[87:80] * 24'h051 + mcu[95:88] * -24'h060 + mcu[103:96] * 24'h060 + mcu[111:104] * -24'h051 + mcu[119:112] * 24'h036 + mcu[127:120] * -24'h013 + mcu[135:128] * -24'h013 + mcu[143:136] * 24'h036 + mcu[151:144] * -24'h051 + mcu[159:152] * 24'h060 + mcu[167:160] * -24'h060 + mcu[175:168] * 24'h051 + mcu[183:176] * -24'h036 + mcu[191:184] * 24'h013 + mcu[199:192] * -24'h02e + mcu[207:200] * 24'h083 + mcu[215:208] * -24'h0c4 + mcu[223:216] * 24'h0e7 + mcu[231:224] * -24'h0e7 + mcu[239:232] * 24'h0c4 + mcu[247:240] * -24'h083 + mcu[255:248] * 24'h02e + mcu[263:256] * -24'h02e + mcu[271:264] * 24'h083 + mcu[279:272] * -24'h0c4 + mcu[287:280] * 24'h0e7 + mcu[295:288] * -24'h0e7 + mcu[303:296] * 24'h0c4 + mcu[311:304] * -24'h083 + mcu[319:312] * 24'h02e + mcu[327:320] * -24'h013 + mcu[335:328] * 24'h036 + mcu[343:336] * -24'h051 + mcu[351:344] * 24'h060 + mcu[359:352] * -24'h060 + mcu[367:360] * 24'h051 + mcu[375:368] * -24'h036 + mcu[383:376] * 24'h013 + mcu[391:384] * 24'h013 + mcu[399:392] * -24'h036 + mcu[407:400] * 24'h051 + mcu[415:408] * -24'h060 + mcu[423:416] * 24'h060 + mcu[431:424] * -24'h051 + mcu[439:432] * 24'h036 + mcu[447:440] * -24'h013 + mcu[455:448] * 24'h02e + mcu[463:456] * -24'h083 + mcu[471:464] * 24'h0c4 + mcu[479:472] * -24'h0e7 + mcu[487:480] * 24'h0e7 + mcu[495:488] * -24'h0c4 + mcu[503:496] * 24'h083 + mcu[511:504] * -24'h02e;
	wire[23:0] cos30_term = mcu[7:0] * 24'h0d4 + mcu[15:8] * 24'h0d4 + mcu[23:16] * 24'h0d4 + mcu[31:24] * 24'h0d4 + mcu[39:32] * 24'h0d4 + mcu[47:40] * 24'h0d4 + mcu[55:48] * 24'h0d4 + mcu[63:56] * 24'h0d4 + mcu[71:64] * -24'h031 + mcu[79:72] * -24'h031 + mcu[87:80] * -24'h031 + mcu[95:88] * -24'h031 + mcu[103:96] * -24'h031 + mcu[111:104] * -24'h031 + mcu[119:112] * -24'h031 + mcu[127:120] * -24'h031 + mcu[135:128] * -24'h0fb + mcu[143:136] * -24'h0fb + mcu[151:144] * -24'h0fb + mcu[159:152] * -24'h0fb + mcu[167:160] * -24'h0fb + mcu[175:168] * -24'h0fb + mcu[183:176] * -24'h0fb + mcu[191:184] * -24'h0fb + mcu[199:192] * -24'h08e + mcu[207:200] * -24'h08e + mcu[215:208] * -24'h08e + mcu[223:216] * -24'h08e + mcu[231:224] * -24'h08e + mcu[239:232] * -24'h08e + mcu[247:240] * -24'h08e + mcu[255:248] * -24'h08e + mcu[263:256] * 24'h08e + mcu[271:264] * 24'h08e + mcu[279:272] * 24'h08e + mcu[287:280] * 24'h08e + mcu[295:288] * 24'h08e + mcu[303:296] * 24'h08e + mcu[311:304] * 24'h08e + mcu[319:312] * 24'h08e + mcu[327:320] * 24'h0fb + mcu[335:328] * 24'h0fb + mcu[343:336] * 24'h0fb + mcu[351:344] * 24'h0fb + mcu[359:352] * 24'h0fb + mcu[367:360] * 24'h0fb + mcu[375:368] * 24'h0fb + mcu[383:376] * 24'h0fb + mcu[391:384] * 24'h031 + mcu[399:392] * 24'h031 + mcu[407:400] * 24'h031 + mcu[415:408] * 24'h031 + mcu[423:416] * 24'h031 + mcu[431:424] * 24'h031 + mcu[439:432] * 24'h031 + mcu[447:440] * 24'h031 + mcu[455:448] * -24'h0d4 + mcu[463:456] * -24'h0d4 + mcu[471:464] * -24'h0d4 + mcu[479:472] * -24'h0d4 + mcu[487:480] * -24'h0d4 + mcu[495:488] * -24'h0d4 + mcu[503:496] * -24'h0d4 + mcu[511:504] * -24'h0d4;
	wire[23:0] cos31_term = mcu[7:0] * 24'h0d0 + mcu[15:8] * 24'h0b0 + mcu[23:16] * 24'h076 + mcu[31:24] * 24'h029 + mcu[39:32] * -24'h029 + mcu[47:40] * -24'h076 + mcu[55:48] * -24'h0b0 + mcu[63:56] * -24'h0d0 + mcu[71:64] * -24'h030 + mcu[79:72] * -24'h029 + mcu[87:80] * -24'h01b + mcu[95:88] * -24'h009 + mcu[103:96] * 24'h009 + mcu[111:104] * 24'h01b + mcu[119:112] * 24'h029 + mcu[127:120] * 24'h030 + mcu[135:128] * -24'h0f6 + mcu[143:136] * -24'h0d0 + mcu[151:144] * -24'h08b + mcu[159:152] * -24'h030 + mcu[167:160] * 24'h030 + mcu[175:168] * 24'h08b + mcu[183:176] * 24'h0d0 + mcu[191:184] * 24'h0f6 + mcu[199:192] * -24'h08b + mcu[207:200] * -24'h076 + mcu[215:208] * -24'h04f + mcu[223:216] * -24'h01b + mcu[231:224] * 24'h01b + mcu[239:232] * 24'h04f + mcu[247:240] * 24'h076 + mcu[255:248] * 24'h08b + mcu[263:256] * 24'h08b + mcu[271:264] * 24'h076 + mcu[279:272] * 24'h04f + mcu[287:280] * 24'h01b + mcu[295:288] * -24'h01b + mcu[303:296] * -24'h04f + mcu[311:304] * -24'h076 + mcu[319:312] * -24'h08b + mcu[327:320] * 24'h0f6 + mcu[335:328] * 24'h0d0 + mcu[343:336] * 24'h08b + mcu[351:344] * 24'h030 + mcu[359:352] * -24'h030 + mcu[367:360] * -24'h08b + mcu[375:368] * -24'h0d0 + mcu[383:376] * -24'h0f6 + mcu[391:384] * 24'h030 + mcu[399:392] * 24'h029 + mcu[407:400] * 24'h01b + mcu[415:408] * 24'h009 + mcu[423:416] * -24'h009 + mcu[431:424] * -24'h01b + mcu[439:432] * -24'h029 + mcu[447:440] * -24'h030 + mcu[455:448] * -24'h0d0 + mcu[463:456] * -24'h0b0 + mcu[471:464] * -24'h076 + mcu[479:472] * -24'h029 + mcu[487:480] * 24'h029 + mcu[495:488] * 24'h076 + mcu[503:496] * 24'h0b0 + mcu[511:504] * 24'h0d0;
	wire[23:0] cos32_term = mcu[7:0] * 24'h0c4 + mcu[15:8] * 24'h051 + mcu[23:16] * -24'h051 + mcu[31:24] * -24'h0c4 + mcu[39:32] * -24'h0c4 + mcu[47:40] * -24'h051 + mcu[55:48] * 24'h051 + mcu[63:56] * 24'h0c4 + mcu[71:64] * -24'h02e + mcu[79:72] * -24'h013 + mcu[87:80] * 24'h013 + mcu[95:88] * 24'h02e + mcu[103:96] * 24'h02e + mcu[111:104] * 24'h013 + mcu[119:112] * -24'h013 + mcu[127:120] * -24'h02e + mcu[135:128] * -24'h0e7 + mcu[143:136] * -24'h060 + mcu[151:144] * 24'h060 + mcu[159:152] * 24'h0e7 + mcu[167:160] * 24'h0e7 + mcu[175:168] * 24'h060 + mcu[183:176] * -24'h060 + mcu[191:184] * -24'h0e7 + mcu[199:192] * -24'h083 + mcu[207:200] * -24'h036 + mcu[215:208] * 24'h036 + mcu[223:216] * 24'h083 + mcu[231:224] * 24'h083 + mcu[239:232] * 24'h036 + mcu[247:240] * -24'h036 + mcu[255:248] * -24'h083 + mcu[263:256] * 24'h083 + mcu[271:264] * 24'h036 + mcu[279:272] * -24'h036 + mcu[287:280] * -24'h083 + mcu[295:288] * -24'h083 + mcu[303:296] * -24'h036 + mcu[311:304] * 24'h036 + mcu[319:312] * 24'h083 + mcu[327:320] * 24'h0e7 + mcu[335:328] * 24'h060 + mcu[343:336] * -24'h060 + mcu[351:344] * -24'h0e7 + mcu[359:352] * -24'h0e7 + mcu[367:360] * -24'h060 + mcu[375:368] * 24'h060 + mcu[383:376] * 24'h0e7 + mcu[391:384] * 24'h02e + mcu[399:392] * 24'h013 + mcu[407:400] * -24'h013 + mcu[415:408] * -24'h02e + mcu[423:416] * -24'h02e + mcu[431:424] * -24'h013 + mcu[439:432] * 24'h013 + mcu[447:440] * 24'h02e + mcu[455:448] * -24'h0c4 + mcu[463:456] * -24'h051 + mcu[471:464] * 24'h051 + mcu[479:472] * 24'h0c4 + mcu[487:480] * 24'h0c4 + mcu[495:488] * 24'h051 + mcu[503:496] * -24'h051 + mcu[511:504] * -24'h0c4;
	wire[23:0] cos33_term = mcu[7:0] * 24'h0b0 + mcu[15:8] * -24'h029 + mcu[23:16] * -24'h0d0 + mcu[31:24] * -24'h076 + mcu[39:32] * 24'h076 + mcu[47:40] * 24'h0d0 + mcu[55:48] * 24'h029 + mcu[63:56] * -24'h0b0 + mcu[71:64] * -24'h029 + mcu[79:72] * 24'h009 + mcu[87:80] * 24'h030 + mcu[95:88] * 24'h01b + mcu[103:96] * -24'h01b + mcu[111:104] * -24'h030 + mcu[119:112] * -24'h009 + mcu[127:120] * 24'h029 + mcu[135:128] * -24'h0d0 + mcu[143:136] * 24'h030 + mcu[151:144] * 24'h0f6 + mcu[159:152] * 24'h08b + mcu[167:160] * -24'h08b + mcu[175:168] * -24'h0f6 + mcu[183:176] * -24'h030 + mcu[191:184] * 24'h0d0 + mcu[199:192] * -24'h076 + mcu[207:200] * 24'h01b + mcu[215:208] * 24'h08b + mcu[223:216] * 24'h04f + mcu[231:224] * -24'h04f + mcu[239:232] * -24'h08b + mcu[247:240] * -24'h01b + mcu[255:248] * 24'h076 + mcu[263:256] * 24'h076 + mcu[271:264] * -24'h01b + mcu[279:272] * -24'h08b + mcu[287:280] * -24'h04f + mcu[295:288] * 24'h04f + mcu[303:296] * 24'h08b + mcu[311:304] * 24'h01b + mcu[319:312] * -24'h076 + mcu[327:320] * 24'h0d0 + mcu[335:328] * -24'h030 + mcu[343:336] * -24'h0f6 + mcu[351:344] * -24'h08b + mcu[359:352] * 24'h08b + mcu[367:360] * 24'h0f6 + mcu[375:368] * 24'h030 + mcu[383:376] * -24'h0d0 + mcu[391:384] * 24'h029 + mcu[399:392] * -24'h009 + mcu[407:400] * -24'h030 + mcu[415:408] * -24'h01b + mcu[423:416] * 24'h01b + mcu[431:424] * 24'h030 + mcu[439:432] * 24'h009 + mcu[447:440] * -24'h029 + mcu[455:448] * -24'h0b0 + mcu[463:456] * 24'h029 + mcu[471:464] * 24'h0d0 + mcu[479:472] * 24'h076 + mcu[487:480] * -24'h076 + mcu[495:488] * -24'h0d0 + mcu[503:496] * -24'h029 + mcu[511:504] * 24'h0b0;
	wire[23:0] cos34_term = mcu[7:0] * 24'h096 + mcu[15:8] * -24'h096 + mcu[23:16] * -24'h096 + mcu[31:24] * 24'h096 + mcu[39:32] * 24'h096 + mcu[47:40] * -24'h096 + mcu[55:48] * -24'h096 + mcu[63:56] * 24'h096 + mcu[71:64] * -24'h023 + mcu[79:72] * 24'h023 + mcu[87:80] * 24'h023 + mcu[95:88] * -24'h023 + mcu[103:96] * -24'h023 + mcu[111:104] * 24'h023 + mcu[119:112] * 24'h023 + mcu[127:120] * -24'h023 + mcu[135:128] * -24'h0b1 + mcu[143:136] * 24'h0b1 + mcu[151:144] * 24'h0b1 + mcu[159:152] * -24'h0b1 + mcu[167:160] * -24'h0b1 + mcu[175:168] * 24'h0b1 + mcu[183:176] * 24'h0b1 + mcu[191:184] * -24'h0b1 + mcu[199:192] * -24'h064 + mcu[207:200] * 24'h064 + mcu[215:208] * 24'h064 + mcu[223:216] * -24'h064 + mcu[231:224] * -24'h064 + mcu[239:232] * 24'h064 + mcu[247:240] * 24'h064 + mcu[255:248] * -24'h064 + mcu[263:256] * 24'h064 + mcu[271:264] * -24'h064 + mcu[279:272] * -24'h064 + mcu[287:280] * 24'h064 + mcu[295:288] * 24'h064 + mcu[303:296] * -24'h064 + mcu[311:304] * -24'h064 + mcu[319:312] * 24'h064 + mcu[327:320] * 24'h0b1 + mcu[335:328] * -24'h0b1 + mcu[343:336] * -24'h0b1 + mcu[351:344] * 24'h0b1 + mcu[359:352] * 24'h0b1 + mcu[367:360] * -24'h0b1 + mcu[375:368] * -24'h0b1 + mcu[383:376] * 24'h0b1 + mcu[391:384] * 24'h023 + mcu[399:392] * -24'h023 + mcu[407:400] * -24'h023 + mcu[415:408] * 24'h023 + mcu[423:416] * 24'h023 + mcu[431:424] * -24'h023 + mcu[439:432] * -24'h023 + mcu[447:440] * 24'h023 + mcu[455:448] * -24'h096 + mcu[463:456] * 24'h096 + mcu[471:464] * 24'h096 + mcu[479:472] * -24'h096 + mcu[487:480] * -24'h096 + mcu[495:488] * 24'h096 + mcu[503:496] * 24'h096 + mcu[511:504] * -24'h096;
	wire[23:0] cos35_term = mcu[7:0] * 24'h076 + mcu[15:8] * -24'h0d0 + mcu[23:16] * 24'h029 + mcu[31:24] * 24'h0b0 + mcu[39:32] * -24'h0b0 + mcu[47:40] * -24'h029 + mcu[55:48] * 24'h0d0 + mcu[63:56] * -24'h076 + mcu[71:64] * -24'h01b + mcu[79:72] * 24'h030 + mcu[87:80] * -24'h009 + mcu[95:88] * -24'h029 + mcu[103:96] * 24'h029 + mcu[111:104] * 24'h009 + mcu[119:112] * -24'h030 + mcu[127:120] * 24'h01b + mcu[135:128] * -24'h08b + mcu[143:136] * 24'h0f6 + mcu[151:144] * -24'h030 + mcu[159:152] * -24'h0d0 + mcu[167:160] * 24'h0d0 + mcu[175:168] * 24'h030 + mcu[183:176] * -24'h0f6 + mcu[191:184] * 24'h08b + mcu[199:192] * -24'h04f + mcu[207:200] * 24'h08b + mcu[215:208] * -24'h01b + mcu[223:216] * -24'h076 + mcu[231:224] * 24'h076 + mcu[239:232] * 24'h01b + mcu[247:240] * -24'h08b + mcu[255:248] * 24'h04f + mcu[263:256] * 24'h04f + mcu[271:264] * -24'h08b + mcu[279:272] * 24'h01b + mcu[287:280] * 24'h076 + mcu[295:288] * -24'h076 + mcu[303:296] * -24'h01b + mcu[311:304] * 24'h08b + mcu[319:312] * -24'h04f + mcu[327:320] * 24'h08b + mcu[335:328] * -24'h0f6 + mcu[343:336] * 24'h030 + mcu[351:344] * 24'h0d0 + mcu[359:352] * -24'h0d0 + mcu[367:360] * -24'h030 + mcu[375:368] * 24'h0f6 + mcu[383:376] * -24'h08b + mcu[391:384] * 24'h01b + mcu[399:392] * -24'h030 + mcu[407:400] * 24'h009 + mcu[415:408] * 24'h029 + mcu[423:416] * -24'h029 + mcu[431:424] * -24'h009 + mcu[439:432] * 24'h030 + mcu[447:440] * -24'h01b + mcu[455:448] * -24'h076 + mcu[463:456] * 24'h0d0 + mcu[471:464] * -24'h029 + mcu[479:472] * -24'h0b0 + mcu[487:480] * 24'h0b0 + mcu[495:488] * 24'h029 + mcu[503:496] * -24'h0d0 + mcu[511:504] * 24'h076;
	wire[23:0] cos36_term = mcu[7:0] * 24'h051 + mcu[15:8] * -24'h0c4 + mcu[23:16] * 24'h0c4 + mcu[31:24] * -24'h051 + mcu[39:32] * -24'h051 + mcu[47:40] * 24'h0c4 + mcu[55:48] * -24'h0c4 + mcu[63:56] * 24'h051 + mcu[71:64] * -24'h013 + mcu[79:72] * 24'h02e + mcu[87:80] * -24'h02e + mcu[95:88] * 24'h013 + mcu[103:96] * 24'h013 + mcu[111:104] * -24'h02e + mcu[119:112] * 24'h02e + mcu[127:120] * -24'h013 + mcu[135:128] * -24'h060 + mcu[143:136] * 24'h0e7 + mcu[151:144] * -24'h0e7 + mcu[159:152] * 24'h060 + mcu[167:160] * 24'h060 + mcu[175:168] * -24'h0e7 + mcu[183:176] * 24'h0e7 + mcu[191:184] * -24'h060 + mcu[199:192] * -24'h036 + mcu[207:200] * 24'h083 + mcu[215:208] * -24'h083 + mcu[223:216] * 24'h036 + mcu[231:224] * 24'h036 + mcu[239:232] * -24'h083 + mcu[247:240] * 24'h083 + mcu[255:248] * -24'h036 + mcu[263:256] * 24'h036 + mcu[271:264] * -24'h083 + mcu[279:272] * 24'h083 + mcu[287:280] * -24'h036 + mcu[295:288] * -24'h036 + mcu[303:296] * 24'h083 + mcu[311:304] * -24'h083 + mcu[319:312] * 24'h036 + mcu[327:320] * 24'h060 + mcu[335:328] * -24'h0e7 + mcu[343:336] * 24'h0e7 + mcu[351:344] * -24'h060 + mcu[359:352] * -24'h060 + mcu[367:360] * 24'h0e7 + mcu[375:368] * -24'h0e7 + mcu[383:376] * 24'h060 + mcu[391:384] * 24'h013 + mcu[399:392] * -24'h02e + mcu[407:400] * 24'h02e + mcu[415:408] * -24'h013 + mcu[423:416] * -24'h013 + mcu[431:424] * 24'h02e + mcu[439:432] * -24'h02e + mcu[447:440] * 24'h013 + mcu[455:448] * -24'h051 + mcu[463:456] * 24'h0c4 + mcu[471:464] * -24'h0c4 + mcu[479:472] * 24'h051 + mcu[487:480] * 24'h051 + mcu[495:488] * -24'h0c4 + mcu[503:496] * 24'h0c4 + mcu[511:504] * -24'h051;
	wire[23:0] cos37_term = mcu[7:0] * 24'h029 + mcu[15:8] * -24'h076 + mcu[23:16] * 24'h0b0 + mcu[31:24] * -24'h0d0 + mcu[39:32] * 24'h0d0 + mcu[47:40] * -24'h0b0 + mcu[55:48] * 24'h076 + mcu[63:56] * -24'h029 + mcu[71:64] * -24'h009 + mcu[79:72] * 24'h01b + mcu[87:80] * -24'h029 + mcu[95:88] * 24'h030 + mcu[103:96] * -24'h030 + mcu[111:104] * 24'h029 + mcu[119:112] * -24'h01b + mcu[127:120] * 24'h009 + mcu[135:128] * -24'h030 + mcu[143:136] * 24'h08b + mcu[151:144] * -24'h0d0 + mcu[159:152] * 24'h0f6 + mcu[167:160] * -24'h0f6 + mcu[175:168] * 24'h0d0 + mcu[183:176] * -24'h08b + mcu[191:184] * 24'h030 + mcu[199:192] * -24'h01b + mcu[207:200] * 24'h04f + mcu[215:208] * -24'h076 + mcu[223:216] * 24'h08b + mcu[231:224] * -24'h08b + mcu[239:232] * 24'h076 + mcu[247:240] * -24'h04f + mcu[255:248] * 24'h01b + mcu[263:256] * 24'h01b + mcu[271:264] * -24'h04f + mcu[279:272] * 24'h076 + mcu[287:280] * -24'h08b + mcu[295:288] * 24'h08b + mcu[303:296] * -24'h076 + mcu[311:304] * 24'h04f + mcu[319:312] * -24'h01b + mcu[327:320] * 24'h030 + mcu[335:328] * -24'h08b + mcu[343:336] * 24'h0d0 + mcu[351:344] * -24'h0f6 + mcu[359:352] * 24'h0f6 + mcu[367:360] * -24'h0d0 + mcu[375:368] * 24'h08b + mcu[383:376] * -24'h030 + mcu[391:384] * 24'h009 + mcu[399:392] * -24'h01b + mcu[407:400] * 24'h029 + mcu[415:408] * -24'h030 + mcu[423:416] * 24'h030 + mcu[431:424] * -24'h029 + mcu[439:432] * 24'h01b + mcu[447:440] * -24'h009 + mcu[455:448] * -24'h029 + mcu[463:456] * 24'h076 + mcu[471:464] * -24'h0b0 + mcu[479:472] * 24'h0d0 + mcu[487:480] * -24'h0d0 + mcu[495:488] * 24'h0b0 + mcu[503:496] * -24'h076 + mcu[511:504] * 24'h029;

	always_comb begin
		dct[15:0] = {cos00_term, 8'b0};
		dct[31:16] = cos01_term;
		dct[47:32] = cos02_term;
		dct[63:48] = cos03_term;
		dct[79:64] = cos04_term;
		dct[95:80] = cos05_term;
		dct[111:96] = cos06_term;
		dct[127:112] = cos07_term;
		dct[143:128] = cos10_term;
		dct[159:144] = cos11_term;
		dct[175:160] = cos12_term;
		dct[191:176] = cos13_term;
		dct[207:192] = cos14_term;
		dct[223:208] = cos15_term;
		dct[239:224] = cos16_term;
		dct[255:240] = cos17_term;
		dct[271:256] = cos20_term;
		dct[287:272] = cos21_term;
		dct[303:288] = cos22_term;
		dct[319:304] = cos23_term;
		dct[335:320] = cos24_term;
		dct[351:336] = cos25_term;
		dct[367:352] = cos26_term;
		dct[383:368] = cos27_term;
		dct[399:384] = cos30_term;
		dct[415:400] = cos31_term;
		dct[431:416] = cos32_term;
		dct[447:432] = cos33_term;
		dct[463:448] = cos34_term;
		dct[479:464] = cos35_term;
		dct[495:480] = cos36_term;
		dct[511:496] = cos37_term;
	end
endmodule
