module dct_quantization(input logic [511:0] mcu, output logic [1023:0] dct);
	wire[47:0] cos00_term = (({8'b0, mcu[7:0], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h100) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h100) >> 8);
	wire[47:0] cos01_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h0fb) >> 8);
	wire[47:0] cos02_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h0ec) >> 8);
	wire[47:0] cos03_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h0d4) >> 8);
	wire[47:0] cos04_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h0b4) >> 8);
	wire[47:0] cos05_term = (({8'b0, mcu[7:0], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h08e) >> 8);
	wire[47:0] cos06_term = (({8'b0, mcu[7:0], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h062) >> 8);
	wire[47:0] cos07_term = (({8'b0, mcu[7:0], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h031) >> 8);
	wire[47:0] cos10_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h0fb) >> 8);
	wire[47:0] cos11_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h0f6) >> 8);
	wire[47:0] cos12_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h0e7) >> 8);
	wire[47:0] cos13_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h0d0) >> 8);
	wire[47:0] cos14_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h0b1) >> 8);
	wire[47:0] cos15_term = (({8'b0, mcu[7:0], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h08b) >> 8);
	wire[47:0] cos16_term = (({8'b0, mcu[7:0], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h060) >> 8);
	wire[47:0] cos17_term = (({8'b0, mcu[7:0], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h030) >> 8);
	wire[47:0] cos20_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h0ec) >> 8);
	wire[47:0] cos21_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h0e7) >> 8);
	wire[47:0] cos22_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h0da) >> 8);
	wire[47:0] cos23_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h0c4) >> 8);
	wire[47:0] cos24_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h0a7) >> 8);
	wire[47:0] cos25_term = (({8'b0, mcu[7:0], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h083) >> 8);
	wire[47:0] cos26_term = (({8'b0, mcu[7:0], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h05a) >> 8);
	wire[47:0] cos27_term = (({8'b0, mcu[7:0], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[71:64], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h02e) >> 8);
	wire[47:0] cos30_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h0d4) >> 8);
	wire[47:0] cos31_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h0d0) >> 8);
	wire[47:0] cos32_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h0c4) >> 8);
	wire[47:0] cos33_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h0b0) >> 8);
	wire[47:0] cos34_term = (({8'b0, mcu[7:0], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h096) >> 8);
	wire[47:0] cos35_term = (({8'b0, mcu[7:0], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h076) >> 8);
	wire[47:0] cos36_term = (({8'b0, mcu[7:0], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h051) >> 8);
	wire[47:0] cos37_term = (({8'b0, mcu[7:0], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h029) >> 8);
	wire[47:0] cos40_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h0b4) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h0b4) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h0b4) >> 8);
	wire[47:0] cos41_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h0b1) >> 8);
	wire[47:0] cos42_term = (({8'b0, mcu[7:0], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h0a7) >> 8);
	wire[47:0] cos43_term = (({8'b0, mcu[7:0], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h096) >> 8);
	wire[47:0] cos44_term = (({8'b0, mcu[7:0], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h080) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h080) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h080) >> 8);
	wire[47:0] cos45_term = (({8'b0, mcu[7:0], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h064) >> 8);
	wire[47:0] cos46_term = (({8'b0, mcu[7:0], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h045) >> 8);
	wire[47:0] cos47_term = (({8'b0, mcu[7:0], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[135:128], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h023) >> 8);
	wire[47:0] cos50_term = (({8'b0, mcu[7:0], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h08e) >> 8);
	wire[47:0] cos51_term = (({8'b0, mcu[7:0], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h08b) >> 8);
	wire[47:0] cos52_term = (({8'b0, mcu[7:0], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h083) >> 8);
	wire[47:0] cos53_term = (({8'b0, mcu[7:0], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h076) >> 8);
	wire[47:0] cos54_term = (({8'b0, mcu[7:0], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h064) >> 8);
	wire[47:0] cos55_term = (({8'b0, mcu[7:0], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h04f) >> 8);
	wire[47:0] cos56_term = (({8'b0, mcu[7:0], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h036) >> 8);
	wire[47:0] cos57_term = (({8'b0, mcu[7:0], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[199:192], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h01b) >> 8);
	wire[47:0] cos60_term = (({8'b0, mcu[7:0], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h062) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h0ec) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h0ec) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h062) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h062) >> 8);
	wire[47:0] cos61_term = (({8'b0, mcu[7:0], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h060) >> 8);
	wire[47:0] cos62_term = (({8'b0, mcu[7:0], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h05a) >> 8);
	wire[47:0] cos63_term = (({8'b0, mcu[7:0], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h051) >> 8);
	wire[47:0] cos64_term = (({8'b0, mcu[7:0], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h0a7) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h0a7) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h045) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h045) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h045) >> 8);
	wire[47:0] cos65_term = (({8'b0, mcu[7:0], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h036) >> 8);
	wire[47:0] cos66_term = (({8'b0, mcu[7:0], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h0da) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h0da) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h025) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h025) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h05a) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h05a) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h025) >> 8);
	wire[47:0] cos67_term = (({8'b0, mcu[7:0], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[263:256], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[327:320], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[391:384], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[455:448], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h013) >> 8);
	wire[47:0] cos70_term = (({8'b0, mcu[7:0], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h031) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h08e) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h0d4) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h0fb) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h0fb) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h0d4) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h08e) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h031) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h031) >> 8);
	wire[47:0] cos71_term = (({8'b0, mcu[7:0], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h030) >> 8);
	wire[47:0] cos72_term = (({8'b0, mcu[7:0], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[15:8], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[79:72], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[143:136], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[207:200], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[271:264], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[335:328], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[399:392], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[463:456], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h02e) >> 8);
	wire[47:0] cos73_term = (({8'b0, mcu[7:0], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h029) >> 8);
	wire[47:0] cos74_term = (({8'b0, mcu[7:0], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[23:16], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[87:80], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[151:144], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[215:208], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[279:272], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h0b1) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h0b1) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[343:336], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h096) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h096) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[407:400], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h064) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h064) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[471:464], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h023) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h023) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h023) >> 8);
	wire[47:0] cos75_term = (({8'b0, mcu[7:0], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[31:24], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[95:88], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[159:152], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[223:216], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[287:280], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[351:344], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[415:408], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[479:472], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h01b) >> 8);
	wire[47:0] cos76_term = (({8'b0, mcu[7:0], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[39:32], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[47:40], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[55:48], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[63:56], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[103:96], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[111:104], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[119:112], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[127:120], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[167:160], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[175:168], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[183:176], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[191:184], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[231:224], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[239:232], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[247:240], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[255:248], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[295:288], 8'b0} * -24'h060) >> 8) + (({8'b0, mcu[303:296], 8'b0} * 24'h0e7) >> 8) + (({8'b0, mcu[311:304], 8'b0} * -24'h0e7) >> 8) + (({8'b0, mcu[319:312], 8'b0} * 24'h060) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[359:352], 8'b0} * 24'h051) >> 8) + (({8'b0, mcu[367:360], 8'b0} * -24'h0c4) >> 8) + (({8'b0, mcu[375:368], 8'b0} * 24'h0c4) >> 8) + (({8'b0, mcu[383:376], 8'b0} * -24'h051) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[423:416], 8'b0} * -24'h036) >> 8) + (({8'b0, mcu[431:424], 8'b0} * 24'h083) >> 8) + (({8'b0, mcu[439:432], 8'b0} * -24'h083) >> 8) + (({8'b0, mcu[447:440], 8'b0} * 24'h036) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h013) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[487:480], 8'b0} * 24'h013) >> 8) + (({8'b0, mcu[495:488], 8'b0} * -24'h02e) >> 8) + (({8'b0, mcu[503:496], 8'b0} * 24'h02e) >> 8) + (({8'b0, mcu[511:504], 8'b0} * -24'h013) >> 8);
	wire[47:0] cos77_term = (({8'b0, mcu[7:0], 8'b0} * 24'h009) >> 8) + (({8'b0, mcu[15:8], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[23:16], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[31:24], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[39:32], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[47:40], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[55:48], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[63:56], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[71:64], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[79:72], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[87:80], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[95:88], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[103:96], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[111:104], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[119:112], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[127:120], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[135:128], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[143:136], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[151:144], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[159:152], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[167:160], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[175:168], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[183:176], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[191:184], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[199:192], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[207:200], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[215:208], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[223:216], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[231:224], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[239:232], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[247:240], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[255:248], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[263:256], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[271:264], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[279:272], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[287:280], 8'b0} * -24'h0f6) >> 8) + (({8'b0, mcu[295:288], 8'b0} * 24'h0f6) >> 8) + (({8'b0, mcu[303:296], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[311:304], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[319:312], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[327:320], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[335:328], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[343:336], 8'b0} * -24'h0b0) >> 8) + (({8'b0, mcu[351:344], 8'b0} * 24'h0d0) >> 8) + (({8'b0, mcu[359:352], 8'b0} * -24'h0d0) >> 8) + (({8'b0, mcu[367:360], 8'b0} * 24'h0b0) >> 8) + (({8'b0, mcu[375:368], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[383:376], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[391:384], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[399:392], 8'b0} * -24'h04f) >> 8) + (({8'b0, mcu[407:400], 8'b0} * 24'h076) >> 8) + (({8'b0, mcu[415:408], 8'b0} * -24'h08b) >> 8) + (({8'b0, mcu[423:416], 8'b0} * 24'h08b) >> 8) + (({8'b0, mcu[431:424], 8'b0} * -24'h076) >> 8) + (({8'b0, mcu[439:432], 8'b0} * 24'h04f) >> 8) + (({8'b0, mcu[447:440], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[455:448], 8'b0} * -24'h009) >> 8) + (({8'b0, mcu[463:456], 8'b0} * 24'h01b) >> 8) + (({8'b0, mcu[471:464], 8'b0} * -24'h029) >> 8) + (({8'b0, mcu[479:472], 8'b0} * 24'h030) >> 8) + (({8'b0, mcu[487:480], 8'b0} * -24'h030) >> 8) + (({8'b0, mcu[495:488], 8'b0} * 24'h029) >> 8) + (({8'b0, mcu[503:496], 8'b0} * -24'h01b) >> 8) + (({8'b0, mcu[511:504], 8'b0} * 24'h009) >> 8);
	
	wire[47:0] cos00_quant = ((cos00_term[23:0] / 24'h10_00) << 8);
	wire[47:0] cos01_quant = ((cos01_term[23:0] / 24'h0B_00) << 8);
	wire[47:0] cos02_quant = ((cos02_term[23:0] / 24'h0A_00) << 8);
	wire[47:0] cos03_quant = ((cos03_term[23:0] / 24'h10_00) << 8);
	wire[47:0] cos04_quant = ((cos04_term[23:0] / 24'h18_00) << 8);
	wire[47:0] cos05_quant = ((cos05_term[23:0] / 24'h28_00) << 8);
	wire[47:0] cos06_quant = ((cos06_term[23:0] / 24'h33_00) << 8);
	wire[47:0] cos07_quant = ((cos07_term[23:0] / 24'h3d_00) << 8);
	wire[47:0] cos10_quant = ((cos10_term[23:0] / 24'h0c_00) << 8);
	wire[47:0] cos11_quant = ((cos11_term[23:0] / 24'h0c_00) << 8);
	wire[47:0] cos12_quant = ((cos12_term[23:0] / 24'h0e_00) << 8);
	wire[47:0] cos13_quant = ((cos13_term[23:0] / 24'h13_00) << 8);
	wire[47:0] cos14_quant = ((cos14_term[23:0] / 24'h1a_00) << 8);
	wire[47:0] cos15_quant = ((cos15_term[23:0] / 24'h3a_00) << 8);
	wire[47:0] cos16_quant = ((cos16_term[23:0] / 24'h3c_00) << 8);
	wire[47:0] cos17_quant = ((cos17_term[23:0] / 24'h37_00) << 8);
	wire[47:0] cos20_quant = ((cos20_term[23:0] / 24'h0e_00) << 8);
	wire[47:0] cos21_quant = ((cos21_term[23:0] / 24'h0d_00) << 8);
	wire[47:0] cos22_quant = ((cos22_term[23:0] / 24'h10_00) << 8);
	wire[47:0] cos23_quant = ((cos23_term[23:0] / 24'h18_00) << 8);
	wire[47:0] cos24_quant = ((cos24_term[23:0] / 24'h28_00) << 8);
	wire[47:0] cos25_quant = ((cos25_term[23:0] / 24'h39_00) << 8);
	wire[47:0] cos26_quant = ((cos26_term[23:0] / 24'h45_00) << 8);
	wire[47:0] cos27_quant = ((cos27_term[23:0] / 24'h38_00) << 8);
	wire[47:0] cos30_quant = ((cos30_term[23:0] / 24'h0e_00) << 8);
	wire[47:0] cos31_quant = ((cos31_term[23:0] / 24'h11_00) << 8);
	wire[47:0] cos32_quant = ((cos32_term[23:0] / 24'h16_00) << 8);
	wire[47:0] cos33_quant = ((cos33_term[23:0] / 24'h1d_00) << 8);
	wire[47:0] cos34_quant = ((cos34_term[23:0] / 24'h33_00) << 8);
	wire[47:0] cos35_quant = ((cos35_term[23:0] / 24'h57_00) << 8);
	wire[47:0] cos36_quant = ((cos36_term[23:0] / 24'h57_00) << 8);
	wire[47:0] cos37_quant = ((cos37_term[23:0] / 24'h3e_00) << 8);
	wire[47:0] cos40_quant = ((cos40_term[23:0] / 24'h12_00) << 8);
	wire[47:0] cos41_quant = ((cos41_term[23:0] / 24'h16_00) << 8);
	wire[47:0] cos42_quant = ((cos42_term[23:0] / 24'h25_00) << 8);
	wire[47:0] cos43_quant = ((cos43_term[23:0] / 24'h38_00) << 8);
	wire[47:0] cos44_quant = ((cos44_term[23:0] / 24'h44_00) << 8);
	wire[47:0] cos45_quant = ((cos45_term[23:0] / 24'h6d_00) << 8);
	wire[47:0] cos46_quant = ((cos46_term[23:0] / 24'h67_00) << 8);
	wire[47:0] cos47_quant = ((cos47_term[23:0] / 24'h4d_00) << 8);
	wire[47:0] cos50_quant = ((cos50_term[23:0] / 24'h18_00) << 8);
	wire[47:0] cos51_quant = ((cos51_term[23:0] / 24'h23_00) << 8);
	wire[47:0] cos52_quant = ((cos52_term[23:0] / 24'h37_00) << 8);
	wire[47:0] cos53_quant = ((cos53_term[23:0] / 24'h40_00) << 8);
	wire[47:0] cos54_quant = ((cos54_term[23:0] / 24'h51_00) << 8);
	wire[47:0] cos55_quant = ((cos55_term[23:0] / 24'h68_00) << 8);
	wire[47:0] cos56_quant = ((cos56_term[23:0] / 24'h71_00) << 8);
	wire[47:0] cos57_quant = ((cos57_term[23:0] / 24'h5c_00) << 8);
	wire[47:0] cos60_quant = ((cos60_term[23:0] / 24'h31_00) << 8);
	wire[47:0] cos61_quant = ((cos61_term[23:0] / 24'h40_00) << 8);
	wire[47:0] cos62_quant = ((cos62_term[23:0] / 24'h4e_00) << 8);
	wire[47:0] cos63_quant = ((cos63_term[23:0] / 24'h57_00) << 8);
	wire[47:0] cos64_quant = ((cos64_term[23:0] / 24'h67_00) << 8);
	wire[47:0] cos65_quant = ((cos65_term[23:0] / 24'h79_00) << 8);
	wire[47:0] cos66_quant = ((cos66_term[23:0] / 24'h78_00) << 8);
	wire[47:0] cos67_quant = ((cos67_term[23:0] / 24'h65_00) << 8);
	wire[47:0] cos70_quant = ((cos70_term[23:0] / 24'h48_00) << 8);
	wire[47:0] cos71_quant = ((cos71_term[23:0] / 24'h5c_00) << 8);
	wire[47:0] cos72_quant = ((cos72_term[23:0] / 24'h5f_00) << 8);
	wire[47:0] cos73_quant = ((cos73_term[23:0] / 24'h62_00) << 8);
	wire[47:0] cos74_quant = ((cos74_term[23:0] / 24'h70_00) << 8);
	wire[47:0] cos75_quant = ((cos75_term[23:0] / 24'h64_00) << 8);
	wire[47:0] cos76_quant = ((cos76_term[23:0] / 24'h67_00) << 8);
	wire[47:0] cos77_quant = ((cos77_term[23:0] / 24'h63_00) << 8);
	always_comb begin
		dct[15:0] = cos00_quant[23:8];
		dct[31:16] = cos01_quant[23:8];
		dct[47:32] = cos02_quant[23:8];
		dct[63:48] = cos03_quant[23:8];
		dct[79:64] = cos04_quant[23:8];
		dct[95:80] = cos05_quant[23:8];
		dct[111:96] = cos06_quant[23:8];
		dct[127:112] = cos07_quant[23:8];
		dct[143:128] = cos10_quant[23:8];
		dct[159:144] = cos11_quant[23:8];
		dct[175:160] = cos12_quant[23:8];
		dct[191:176] = cos13_quant[23:8];
		dct[207:192] = cos14_quant[23:8];
		dct[223:208] = cos15_quant[23:8];
		dct[239:224] = cos16_quant[23:8];
		dct[255:240] = cos17_quant[23:8];
		dct[271:256] = cos20_quant[23:8];
		dct[287:272] = cos21_quant[23:8];
		dct[303:288] = cos22_quant[23:8];
		dct[319:304] = cos23_quant[23:8];
		dct[335:320] = cos24_quant[23:8];
		dct[351:336] = cos25_quant[23:8];
		dct[367:352] = cos26_quant[23:8];
		dct[383:368] = cos27_quant[23:8];
		dct[399:384] = cos30_quant[23:8];
		dct[415:400] = cos31_quant[23:8];
		dct[431:416] = cos32_quant[23:8];
		dct[447:432] = cos33_quant[23:8];
		dct[463:448] = cos34_quant[23:8];
		dct[479:464] = cos35_quant[23:8];
		dct[495:480] = cos36_quant[23:8];
		dct[511:496] = cos37_quant[23:8];
		dct[527:512] = cos40_quant[23:8];
		dct[543:528] = cos41_quant[23:8];
		dct[559:544] = cos42_quant[23:8];
		dct[575:560] = cos43_quant[23:8];
		dct[591:576] = cos44_quant[23:8];
		dct[607:592] = cos45_quant[23:8];
		dct[623:608] = cos46_quant[23:8];
		dct[639:624] = cos47_quant[23:8];
		dct[655:640] = cos50_quant[23:8];
		dct[671:656] = cos51_quant[23:8];
		dct[687:672] = cos52_quant[23:8];
		dct[703:688] = cos53_quant[23:8];
		dct[719:704] = cos54_quant[23:8];
		dct[735:720] = cos55_quant[23:8];
		dct[751:736] = cos56_quant[23:8];
		dct[767:752] = cos57_quant[23:8];
		dct[783:768] = cos60_quant[23:8];
		dct[799:784] = cos61_quant[23:8];
		dct[815:800] = cos62_quant[23:8];
		dct[831:816] = cos63_quant[23:8];
		dct[847:832] = cos64_quant[23:8];
		dct[863:848] = cos65_quant[23:8];
		dct[879:864] = cos66_quant[23:8];
		dct[895:880] = cos67_quant[23:8];
		dct[911:896] = cos70_quant[23:8];
		dct[927:912] = cos71_quant[23:8];
		dct[943:928] = cos72_quant[23:8];
		dct[959:944] = cos73_quant[23:8];
		dct[975:960] = cos74_quant[23:8];
		dct[991:976] = cos75_quant[23:8];
		dct[1007:992] = cos76_quant[23:8];
		dct[1023:1008] = cos77_quant[23:8];
	end
endmodule