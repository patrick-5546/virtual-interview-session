module dct_quantization(input logic [511:0] mcu, output logic [1023:0] dct);
	wire[15:0] cos00_term = mcu[7:0] + mcu[15:8] + mcu[23:16] + mcu[31:24] + mcu[39:32] + mcu[47:40] + mcu[55:48] + mcu[63:56] + mcu[71:64] + mcu[79:72] + mcu[87:80] + mcu[95:88] + mcu[103:96] + mcu[111:104] + mcu[119:112] + mcu[127:120] + mcu[135:128] + mcu[143:136] + mcu[151:144] + mcu[159:152] + mcu[167:160] + mcu[175:168] + mcu[183:176] + mcu[191:184] + mcu[199:192] + mcu[207:200] + mcu[215:208] + mcu[223:216] + mcu[231:224] + mcu[239:232] + mcu[247:240] + mcu[255:248] + mcu[263:256] + mcu[271:264] + mcu[279:272] + mcu[287:280] + mcu[295:288] + mcu[303:296] + mcu[311:304] + mcu[319:312] + mcu[327:320] + mcu[335:328] + mcu[343:336] + mcu[351:344] + mcu[359:352] + mcu[367:360] + mcu[375:368] + mcu[383:376] + mcu[391:384] + mcu[399:392] + mcu[407:400] + mcu[415:408] + mcu[423:416] + mcu[431:424] + mcu[439:432] + mcu[447:440] + mcu[455:448] + mcu[463:456] + mcu[471:464] + mcu[479:472] + mcu[487:480] + mcu[495:488] + mcu[503:496] + mcu[511:504];
	wire[23:0] cos01_term = mcu[7:0] * 24'h0fb + mcu[15:8] * 24'h0d4 + mcu[23:16] * 24'h08e + mcu[31:24] * 24'h031 + mcu[39:32] * -24'h031 + mcu[47:40] * -24'h08e + mcu[55:48] * -24'h0d4 + mcu[63:56] * -24'h0fb + mcu[71:64] * 24'h0fb + mcu[79:72] * 24'h0d4 + mcu[87:80] * 24'h08e + mcu[95:88] * 24'h031 + mcu[103:96] * -24'h031 + mcu[111:104] * -24'h08e + mcu[119:112] * -24'h0d4 + mcu[127:120] * -24'h0fb + mcu[135:128] * 24'h0fb + mcu[143:136] * 24'h0d4 + mcu[151:144] * 24'h08e + mcu[159:152] * 24'h031 + mcu[167:160] * -24'h031 + mcu[175:168] * -24'h08e + mcu[183:176] * -24'h0d4 + mcu[191:184] * -24'h0fb + mcu[199:192] * 24'h0fb + mcu[207:200] * 24'h0d4 + mcu[215:208] * 24'h08e + mcu[223:216] * 24'h031 + mcu[231:224] * -24'h031 + mcu[239:232] * -24'h08e + mcu[247:240] * -24'h0d4 + mcu[255:248] * -24'h0fb + mcu[263:256] * 24'h0fb + mcu[271:264] * 24'h0d4 + mcu[279:272] * 24'h08e + mcu[287:280] * 24'h031 + mcu[295:288] * -24'h031 + mcu[303:296] * -24'h08e + mcu[311:304] * -24'h0d4 + mcu[319:312] * -24'h0fb + mcu[327:320] * 24'h0fb + mcu[335:328] * 24'h0d4 + mcu[343:336] * 24'h08e + mcu[351:344] * 24'h031 + mcu[359:352] * -24'h031 + mcu[367:360] * -24'h08e + mcu[375:368] * -24'h0d4 + mcu[383:376] * -24'h0fb + mcu[391:384] * 24'h0fb + mcu[399:392] * 24'h0d4 + mcu[407:400] * 24'h08e + mcu[415:408] * 24'h031 + mcu[423:416] * -24'h031 + mcu[431:424] * -24'h08e + mcu[439:432] * -24'h0d4 + mcu[447:440] * -24'h0fb + mcu[455:448] * 24'h0fb + mcu[463:456] * 24'h0d4 + mcu[471:464] * 24'h08e + mcu[479:472] * 24'h031 + mcu[487:480] * -24'h031 + mcu[495:488] * -24'h08e + mcu[503:496] * -24'h0d4 + mcu[511:504] * -24'h0fb;
	wire[47:0] cos02_term = (({mcu[7:0], 8'b0} * 24'h0ec)) + (({mcu[15:8], 8'b0} * 24'h062)) + (({mcu[23:16], 8'b0} * -24'h062)) + (({mcu[31:24], 8'b0} * -24'h0ec)) + (({mcu[39:32], 8'b0} * -24'h0ec)) + (({mcu[47:40], 8'b0} * -24'h062)) + (({mcu[55:48], 8'b0} * 24'h062)) + (({mcu[63:56], 8'b0} * 24'h0ec)) + (({mcu[71:64], 8'b0} * 24'h0ec)) + (({mcu[79:72], 8'b0} * 24'h062)) + (({mcu[87:80], 8'b0} * -24'h062)) + (({mcu[95:88], 8'b0} * -24'h0ec)) + (({mcu[103:96], 8'b0} * -24'h0ec)) + (({mcu[111:104], 8'b0} * -24'h062)) + (({mcu[119:112], 8'b0} * 24'h062)) + (({mcu[127:120], 8'b0} * 24'h0ec)) + (({mcu[135:128], 8'b0} * 24'h0ec)) + (({mcu[143:136], 8'b0} * 24'h062)) + (({mcu[151:144], 8'b0} * -24'h062)) + (({mcu[159:152], 8'b0} * -24'h0ec)) + (({mcu[167:160], 8'b0} * -24'h0ec)) + (({mcu[175:168], 8'b0} * -24'h062)) + (({mcu[183:176], 8'b0} * 24'h062)) + (({mcu[191:184], 8'b0} * 24'h0ec)) + (({mcu[199:192], 8'b0} * 24'h0ec)) + (({mcu[207:200], 8'b0} * 24'h062)) + (({mcu[215:208], 8'b0} * -24'h062)) + (({mcu[223:216], 8'b0} * -24'h0ec)) + (({mcu[231:224], 8'b0} * -24'h0ec)) + (({mcu[239:232], 8'b0} * -24'h062)) + (({mcu[247:240], 8'b0} * 24'h062)) + (({mcu[255:248], 8'b0} * 24'h0ec)) + (({mcu[263:256], 8'b0} * 24'h0ec)) + (({mcu[271:264], 8'b0} * 24'h062)) + (({mcu[279:272], 8'b0} * -24'h062)) + (({mcu[287:280], 8'b0} * -24'h0ec)) + (({mcu[295:288], 8'b0} * -24'h0ec)) + (({mcu[303:296], 8'b0} * -24'h062)) + (({mcu[311:304], 8'b0} * 24'h062)) + (({mcu[319:312], 8'b0} * 24'h0ec)) + (({mcu[327:320], 8'b0} * 24'h0ec)) + (({mcu[335:328], 8'b0} * 24'h062)) + (({mcu[343:336], 8'b0} * -24'h062)) + (({mcu[351:344], 8'b0} * -24'h0ec)) + (({mcu[359:352], 8'b0} * -24'h0ec)) + (({mcu[367:360], 8'b0} * -24'h062)) + (({mcu[375:368], 8'b0} * 24'h062)) + (({mcu[383:376], 8'b0} * 24'h0ec)) + (({mcu[391:384], 8'b0} * 24'h0ec)) + (({mcu[399:392], 8'b0} * 24'h062)) + (({mcu[407:400], 8'b0} * -24'h062)) + (({mcu[415:408], 8'b0} * -24'h0ec)) + (({mcu[423:416], 8'b0} * -24'h0ec)) + (({mcu[431:424], 8'b0} * -24'h062)) + (({mcu[439:432], 8'b0} * 24'h062)) + (({mcu[447:440], 8'b0} * 24'h0ec)) + (({mcu[455:448], 8'b0} * 24'h0ec)) + (({mcu[463:456], 8'b0} * 24'h062)) + (({mcu[471:464], 8'b0} * -24'h062)) + (({mcu[479:472], 8'b0} * -24'h0ec)) + (({mcu[487:480], 8'b0} * -24'h0ec)) + (({mcu[495:488], 8'b0} * -24'h062)) + (({mcu[503:496], 8'b0} * 24'h062)) + (({mcu[511:504], 8'b0} * 24'h0ec));
	wire[47:0] cos03_term = (({mcu[7:0], 8'b0} * 24'h0d4)) + (({mcu[15:8], 8'b0} * -24'h031)) + (({mcu[23:16], 8'b0} * -24'h0fb)) + (({mcu[31:24], 8'b0} * -24'h08e)) + (({mcu[39:32], 8'b0} * 24'h08e)) + (({mcu[47:40], 8'b0} * 24'h0fb)) + (({mcu[55:48], 8'b0} * 24'h031)) + (({mcu[63:56], 8'b0} * -24'h0d4)) + (({mcu[71:64], 8'b0} * 24'h0d4)) + (({mcu[79:72], 8'b0} * -24'h031)) + (({mcu[87:80], 8'b0} * -24'h0fb)) + (({mcu[95:88], 8'b0} * -24'h08e)) + (({mcu[103:96], 8'b0} * 24'h08e)) + (({mcu[111:104], 8'b0} * 24'h0fb)) + (({mcu[119:112], 8'b0} * 24'h031)) + (({mcu[127:120], 8'b0} * -24'h0d4)) + (({mcu[135:128], 8'b0} * 24'h0d4)) + (({mcu[143:136], 8'b0} * -24'h031)) + (({mcu[151:144], 8'b0} * -24'h0fb)) + (({mcu[159:152], 8'b0} * -24'h08e)) + (({mcu[167:160], 8'b0} * 24'h08e)) + (({mcu[175:168], 8'b0} * 24'h0fb)) + (({mcu[183:176], 8'b0} * 24'h031)) + (({mcu[191:184], 8'b0} * -24'h0d4)) + (({mcu[199:192], 8'b0} * 24'h0d4)) + (({mcu[207:200], 8'b0} * -24'h031)) + (({mcu[215:208], 8'b0} * -24'h0fb)) + (({mcu[223:216], 8'b0} * -24'h08e)) + (({mcu[231:224], 8'b0} * 24'h08e)) + (({mcu[239:232], 8'b0} * 24'h0fb)) + (({mcu[247:240], 8'b0} * 24'h031)) + (({mcu[255:248], 8'b0} * -24'h0d4)) + (({mcu[263:256], 8'b0} * 24'h0d4)) + (({mcu[271:264], 8'b0} * -24'h031)) + (({mcu[279:272], 8'b0} * -24'h0fb)) + (({mcu[287:280], 8'b0} * -24'h08e)) + (({mcu[295:288], 8'b0} * 24'h08e)) + (({mcu[303:296], 8'b0} * 24'h0fb)) + (({mcu[311:304], 8'b0} * 24'h031)) + (({mcu[319:312], 8'b0} * -24'h0d4)) + (({mcu[327:320], 8'b0} * 24'h0d4)) + (({mcu[335:328], 8'b0} * -24'h031)) + (({mcu[343:336], 8'b0} * -24'h0fb)) + (({mcu[351:344], 8'b0} * -24'h08e)) + (({mcu[359:352], 8'b0} * 24'h08e)) + (({mcu[367:360], 8'b0} * 24'h0fb)) + (({mcu[375:368], 8'b0} * 24'h031)) + (({mcu[383:376], 8'b0} * -24'h0d4)) + (({mcu[391:384], 8'b0} * 24'h0d4)) + (({mcu[399:392], 8'b0} * -24'h031)) + (({mcu[407:400], 8'b0} * -24'h0fb)) + (({mcu[415:408], 8'b0} * -24'h08e)) + (({mcu[423:416], 8'b0} * 24'h08e)) + (({mcu[431:424], 8'b0} * 24'h0fb)) + (({mcu[439:432], 8'b0} * 24'h031)) + (({mcu[447:440], 8'b0} * -24'h0d4)) + (({mcu[455:448], 8'b0} * 24'h0d4)) + (({mcu[463:456], 8'b0} * -24'h031)) + (({mcu[471:464], 8'b0} * -24'h0fb)) + (({mcu[479:472], 8'b0} * -24'h08e)) + (({mcu[487:480], 8'b0} * 24'h08e)) + (({mcu[495:488], 8'b0} * 24'h0fb)) + (({mcu[503:496], 8'b0} * 24'h031)) + (({mcu[511:504], 8'b0} * -24'h0d4));
	wire[47:0] cos04_term = (({mcu[7:0], 8'b0} * 24'h0b4)) + (({mcu[15:8], 8'b0} * -24'h0b4)) + (({mcu[23:16], 8'b0} * -24'h0b4)) + (({mcu[31:24], 8'b0} * 24'h0b4)) + (({mcu[39:32], 8'b0} * 24'h0b4)) + (({mcu[47:40], 8'b0} * -24'h0b4)) + (({mcu[55:48], 8'b0} * -24'h0b4)) + (({mcu[63:56], 8'b0} * 24'h0b4)) + (({mcu[71:64], 8'b0} * 24'h0b4)) + (({mcu[79:72], 8'b0} * -24'h0b4)) + (({mcu[87:80], 8'b0} * -24'h0b4)) + (({mcu[95:88], 8'b0} * 24'h0b4)) + (({mcu[103:96], 8'b0} * 24'h0b4)) + (({mcu[111:104], 8'b0} * -24'h0b4)) + (({mcu[119:112], 8'b0} * -24'h0b4)) + (({mcu[127:120], 8'b0} * 24'h0b4)) + (({mcu[135:128], 8'b0} * 24'h0b4)) + (({mcu[143:136], 8'b0} * -24'h0b4)) + (({mcu[151:144], 8'b0} * -24'h0b4)) + (({mcu[159:152], 8'b0} * 24'h0b4)) + (({mcu[167:160], 8'b0} * 24'h0b4)) + (({mcu[175:168], 8'b0} * -24'h0b4)) + (({mcu[183:176], 8'b0} * -24'h0b4)) + (({mcu[191:184], 8'b0} * 24'h0b4)) + (({mcu[199:192], 8'b0} * 24'h0b4)) + (({mcu[207:200], 8'b0} * -24'h0b4)) + (({mcu[215:208], 8'b0} * -24'h0b4)) + (({mcu[223:216], 8'b0} * 24'h0b4)) + (({mcu[231:224], 8'b0} * 24'h0b4)) + (({mcu[239:232], 8'b0} * -24'h0b4)) + (({mcu[247:240], 8'b0} * -24'h0b4)) + (({mcu[255:248], 8'b0} * 24'h0b4)) + (({mcu[263:256], 8'b0} * 24'h0b4)) + (({mcu[271:264], 8'b0} * -24'h0b4)) + (({mcu[279:272], 8'b0} * -24'h0b4)) + (({mcu[287:280], 8'b0} * 24'h0b4)) + (({mcu[295:288], 8'b0} * 24'h0b4)) + (({mcu[303:296], 8'b0} * -24'h0b4)) + (({mcu[311:304], 8'b0} * -24'h0b4)) + (({mcu[319:312], 8'b0} * 24'h0b4)) + (({mcu[327:320], 8'b0} * 24'h0b4)) + (({mcu[335:328], 8'b0} * -24'h0b4)) + (({mcu[343:336], 8'b0} * -24'h0b4)) + (({mcu[351:344], 8'b0} * 24'h0b4)) + (({mcu[359:352], 8'b0} * 24'h0b4)) + (({mcu[367:360], 8'b0} * -24'h0b4)) + (({mcu[375:368], 8'b0} * -24'h0b4)) + (({mcu[383:376], 8'b0} * 24'h0b4)) + (({mcu[391:384], 8'b0} * 24'h0b4)) + (({mcu[399:392], 8'b0} * -24'h0b4)) + (({mcu[407:400], 8'b0} * -24'h0b4)) + (({mcu[415:408], 8'b0} * 24'h0b4)) + (({mcu[423:416], 8'b0} * 24'h0b4)) + (({mcu[431:424], 8'b0} * -24'h0b4)) + (({mcu[439:432], 8'b0} * -24'h0b4)) + (({mcu[447:440], 8'b0} * 24'h0b4)) + (({mcu[455:448], 8'b0} * 24'h0b4)) + (({mcu[463:456], 8'b0} * -24'h0b4)) + (({mcu[471:464], 8'b0} * -24'h0b4)) + (({mcu[479:472], 8'b0} * 24'h0b4)) + (({mcu[487:480], 8'b0} * 24'h0b4)) + (({mcu[495:488], 8'b0} * -24'h0b4)) + (({mcu[503:496], 8'b0} * -24'h0b4)) + (({mcu[511:504], 8'b0} * 24'h0b4));
	wire[47:0] cos05_term = (({mcu[7:0], 8'b0} * 24'h08e)) + (({mcu[15:8], 8'b0} * -24'h0fb)) + (({mcu[23:16], 8'b0} * 24'h031)) + (({mcu[31:24], 8'b0} * 24'h0d4)) + (({mcu[39:32], 8'b0} * -24'h0d4)) + (({mcu[47:40], 8'b0} * -24'h031)) + (({mcu[55:48], 8'b0} * 24'h0fb)) + (({mcu[63:56], 8'b0} * -24'h08e)) + (({mcu[71:64], 8'b0} * 24'h08e)) + (({mcu[79:72], 8'b0} * -24'h0fb)) + (({mcu[87:80], 8'b0} * 24'h031)) + (({mcu[95:88], 8'b0} * 24'h0d4)) + (({mcu[103:96], 8'b0} * -24'h0d4)) + (({mcu[111:104], 8'b0} * -24'h031)) + (({mcu[119:112], 8'b0} * 24'h0fb)) + (({mcu[127:120], 8'b0} * -24'h08e)) + (({mcu[135:128], 8'b0} * 24'h08e)) + (({mcu[143:136], 8'b0} * -24'h0fb)) + (({mcu[151:144], 8'b0} * 24'h031)) + (({mcu[159:152], 8'b0} * 24'h0d4)) + (({mcu[167:160], 8'b0} * -24'h0d4)) + (({mcu[175:168], 8'b0} * -24'h031)) + (({mcu[183:176], 8'b0} * 24'h0fb)) + (({mcu[191:184], 8'b0} * -24'h08e)) + (({mcu[199:192], 8'b0} * 24'h08e)) + (({mcu[207:200], 8'b0} * -24'h0fb)) + (({mcu[215:208], 8'b0} * 24'h031)) + (({mcu[223:216], 8'b0} * 24'h0d4)) + (({mcu[231:224], 8'b0} * -24'h0d4)) + (({mcu[239:232], 8'b0} * -24'h031)) + (({mcu[247:240], 8'b0} * 24'h0fb)) + (({mcu[255:248], 8'b0} * -24'h08e)) + (({mcu[263:256], 8'b0} * 24'h08e)) + (({mcu[271:264], 8'b0} * -24'h0fb)) + (({mcu[279:272], 8'b0} * 24'h031)) + (({mcu[287:280], 8'b0} * 24'h0d4)) + (({mcu[295:288], 8'b0} * -24'h0d4)) + (({mcu[303:296], 8'b0} * -24'h031)) + (({mcu[311:304], 8'b0} * 24'h0fb)) + (({mcu[319:312], 8'b0} * -24'h08e)) + (({mcu[327:320], 8'b0} * 24'h08e)) + (({mcu[335:328], 8'b0} * -24'h0fb)) + (({mcu[343:336], 8'b0} * 24'h031)) + (({mcu[351:344], 8'b0} * 24'h0d4)) + (({mcu[359:352], 8'b0} * -24'h0d4)) + (({mcu[367:360], 8'b0} * -24'h031)) + (({mcu[375:368], 8'b0} * 24'h0fb)) + (({mcu[383:376], 8'b0} * -24'h08e)) + (({mcu[391:384], 8'b0} * 24'h08e)) + (({mcu[399:392], 8'b0} * -24'h0fb)) + (({mcu[407:400], 8'b0} * 24'h031)) + (({mcu[415:408], 8'b0} * 24'h0d4)) + (({mcu[423:416], 8'b0} * -24'h0d4)) + (({mcu[431:424], 8'b0} * -24'h031)) + (({mcu[439:432], 8'b0} * 24'h0fb)) + (({mcu[447:440], 8'b0} * -24'h08e)) + (({mcu[455:448], 8'b0} * 24'h08e)) + (({mcu[463:456], 8'b0} * -24'h0fb)) + (({mcu[471:464], 8'b0} * 24'h031)) + (({mcu[479:472], 8'b0} * 24'h0d4)) + (({mcu[487:480], 8'b0} * -24'h0d4)) + (({mcu[495:488], 8'b0} * -24'h031)) + (({mcu[503:496], 8'b0} * 24'h0fb)) + (({mcu[511:504], 8'b0} * -24'h08e));
	wire[47:0] cos06_term = (({mcu[7:0], 8'b0} * 24'h062)) + (({mcu[15:8], 8'b0} * -24'h0ec)) + (({mcu[23:16], 8'b0} * 24'h0ec)) + (({mcu[31:24], 8'b0} * -24'h062)) + (({mcu[39:32], 8'b0} * -24'h062)) + (({mcu[47:40], 8'b0} * 24'h0ec)) + (({mcu[55:48], 8'b0} * -24'h0ec)) + (({mcu[63:56], 8'b0} * 24'h062)) + (({mcu[71:64], 8'b0} * 24'h062)) + (({mcu[79:72], 8'b0} * -24'h0ec)) + (({mcu[87:80], 8'b0} * 24'h0ec)) + (({mcu[95:88], 8'b0} * -24'h062)) + (({mcu[103:96], 8'b0} * -24'h062)) + (({mcu[111:104], 8'b0} * 24'h0ec)) + (({mcu[119:112], 8'b0} * -24'h0ec)) + (({mcu[127:120], 8'b0} * 24'h062)) + (({mcu[135:128], 8'b0} * 24'h062)) + (({mcu[143:136], 8'b0} * -24'h0ec)) + (({mcu[151:144], 8'b0} * 24'h0ec)) + (({mcu[159:152], 8'b0} * -24'h062)) + (({mcu[167:160], 8'b0} * -24'h062)) + (({mcu[175:168], 8'b0} * 24'h0ec)) + (({mcu[183:176], 8'b0} * -24'h0ec)) + (({mcu[191:184], 8'b0} * 24'h062)) + (({mcu[199:192], 8'b0} * 24'h062)) + (({mcu[207:200], 8'b0} * -24'h0ec)) + (({mcu[215:208], 8'b0} * 24'h0ec)) + (({mcu[223:216], 8'b0} * -24'h062)) + (({mcu[231:224], 8'b0} * -24'h062)) + (({mcu[239:232], 8'b0} * 24'h0ec)) + (({mcu[247:240], 8'b0} * -24'h0ec)) + (({mcu[255:248], 8'b0} * 24'h062)) + (({mcu[263:256], 8'b0} * 24'h062)) + (({mcu[271:264], 8'b0} * -24'h0ec)) + (({mcu[279:272], 8'b0} * 24'h0ec)) + (({mcu[287:280], 8'b0} * -24'h062)) + (({mcu[295:288], 8'b0} * -24'h062)) + (({mcu[303:296], 8'b0} * 24'h0ec)) + (({mcu[311:304], 8'b0} * -24'h0ec)) + (({mcu[319:312], 8'b0} * 24'h062)) + (({mcu[327:320], 8'b0} * 24'h062)) + (({mcu[335:328], 8'b0} * -24'h0ec)) + (({mcu[343:336], 8'b0} * 24'h0ec)) + (({mcu[351:344], 8'b0} * -24'h062)) + (({mcu[359:352], 8'b0} * -24'h062)) + (({mcu[367:360], 8'b0} * 24'h0ec)) + (({mcu[375:368], 8'b0} * -24'h0ec)) + (({mcu[383:376], 8'b0} * 24'h062)) + (({mcu[391:384], 8'b0} * 24'h062)) + (({mcu[399:392], 8'b0} * -24'h0ec)) + (({mcu[407:400], 8'b0} * 24'h0ec)) + (({mcu[415:408], 8'b0} * -24'h062)) + (({mcu[423:416], 8'b0} * -24'h062)) + (({mcu[431:424], 8'b0} * 24'h0ec)) + (({mcu[439:432], 8'b0} * -24'h0ec)) + (({mcu[447:440], 8'b0} * 24'h062)) + (({mcu[455:448], 8'b0} * 24'h062)) + (({mcu[463:456], 8'b0} * -24'h0ec)) + (({mcu[471:464], 8'b0} * 24'h0ec)) + (({mcu[479:472], 8'b0} * -24'h062)) + (({mcu[487:480], 8'b0} * -24'h062)) + (({mcu[495:488], 8'b0} * 24'h0ec)) + (({mcu[503:496], 8'b0} * -24'h0ec)) + (({mcu[511:504], 8'b0} * 24'h062));
	wire[47:0] cos07_term = (({mcu[7:0], 8'b0} * 24'h031)) + (({mcu[15:8], 8'b0} * -24'h08e)) + (({mcu[23:16], 8'b0} * 24'h0d4)) + (({mcu[31:24], 8'b0} * -24'h0fb)) + (({mcu[39:32], 8'b0} * 24'h0fb)) + (({mcu[47:40], 8'b0} * -24'h0d4)) + (({mcu[55:48], 8'b0} * 24'h08e)) + (({mcu[63:56], 8'b0} * -24'h031)) + (({mcu[71:64], 8'b0} * 24'h031)) + (({mcu[79:72], 8'b0} * -24'h08e)) + (({mcu[87:80], 8'b0} * 24'h0d4)) + (({mcu[95:88], 8'b0} * -24'h0fb)) + (({mcu[103:96], 8'b0} * 24'h0fb)) + (({mcu[111:104], 8'b0} * -24'h0d4)) + (({mcu[119:112], 8'b0} * 24'h08e)) + (({mcu[127:120], 8'b0} * -24'h031)) + (({mcu[135:128], 8'b0} * 24'h031)) + (({mcu[143:136], 8'b0} * -24'h08e)) + (({mcu[151:144], 8'b0} * 24'h0d4)) + (({mcu[159:152], 8'b0} * -24'h0fb)) + (({mcu[167:160], 8'b0} * 24'h0fb)) + (({mcu[175:168], 8'b0} * -24'h0d4)) + (({mcu[183:176], 8'b0} * 24'h08e)) + (({mcu[191:184], 8'b0} * -24'h031)) + (({mcu[199:192], 8'b0} * 24'h031)) + (({mcu[207:200], 8'b0} * -24'h08e)) + (({mcu[215:208], 8'b0} * 24'h0d4)) + (({mcu[223:216], 8'b0} * -24'h0fb)) + (({mcu[231:224], 8'b0} * 24'h0fb)) + (({mcu[239:232], 8'b0} * -24'h0d4)) + (({mcu[247:240], 8'b0} * 24'h08e)) + (({mcu[255:248], 8'b0} * -24'h031)) + (({mcu[263:256], 8'b0} * 24'h031)) + (({mcu[271:264], 8'b0} * -24'h08e)) + (({mcu[279:272], 8'b0} * 24'h0d4)) + (({mcu[287:280], 8'b0} * -24'h0fb)) + (({mcu[295:288], 8'b0} * 24'h0fb)) + (({mcu[303:296], 8'b0} * -24'h0d4)) + (({mcu[311:304], 8'b0} * 24'h08e)) + (({mcu[319:312], 8'b0} * -24'h031)) + (({mcu[327:320], 8'b0} * 24'h031)) + (({mcu[335:328], 8'b0} * -24'h08e)) + (({mcu[343:336], 8'b0} * 24'h0d4)) + (({mcu[351:344], 8'b0} * -24'h0fb)) + (({mcu[359:352], 8'b0} * 24'h0fb)) + (({mcu[367:360], 8'b0} * -24'h0d4)) + (({mcu[375:368], 8'b0} * 24'h08e)) + (({mcu[383:376], 8'b0} * -24'h031)) + (({mcu[391:384], 8'b0} * 24'h031)) + (({mcu[399:392], 8'b0} * -24'h08e)) + (({mcu[407:400], 8'b0} * 24'h0d4)) + (({mcu[415:408], 8'b0} * -24'h0fb)) + (({mcu[423:416], 8'b0} * 24'h0fb)) + (({mcu[431:424], 8'b0} * -24'h0d4)) + (({mcu[439:432], 8'b0} * 24'h08e)) + (({mcu[447:440], 8'b0} * -24'h031)) + (({mcu[455:448], 8'b0} * 24'h031)) + (({mcu[463:456], 8'b0} * -24'h08e)) + (({mcu[471:464], 8'b0} * 24'h0d4)) + (({mcu[479:472], 8'b0} * -24'h0fb)) + (({mcu[487:480], 8'b0} * 24'h0fb)) + (({mcu[495:488], 8'b0} * -24'h0d4)) + (({mcu[503:496], 8'b0} * 24'h08e)) + (({mcu[511:504], 8'b0} * -24'h031));
	wire[47:0] cos10_term = (({mcu[7:0], 8'b0} * 24'h0fb)) + (({mcu[15:8], 8'b0} * 24'h0fb)) + (({mcu[23:16], 8'b0} * 24'h0fb)) + (({mcu[31:24], 8'b0} * 24'h0fb)) + (({mcu[39:32], 8'b0} * 24'h0fb)) + (({mcu[47:40], 8'b0} * 24'h0fb)) + (({mcu[55:48], 8'b0} * 24'h0fb)) + (({mcu[63:56], 8'b0} * 24'h0fb)) + (({mcu[71:64], 8'b0} * 24'h0d4)) + (({mcu[79:72], 8'b0} * 24'h0d4)) + (({mcu[87:80], 8'b0} * 24'h0d4)) + (({mcu[95:88], 8'b0} * 24'h0d4)) + (({mcu[103:96], 8'b0} * 24'h0d4)) + (({mcu[111:104], 8'b0} * 24'h0d4)) + (({mcu[119:112], 8'b0} * 24'h0d4)) + (({mcu[127:120], 8'b0} * 24'h0d4)) + (({mcu[135:128], 8'b0} * 24'h08e)) + (({mcu[143:136], 8'b0} * 24'h08e)) + (({mcu[151:144], 8'b0} * 24'h08e)) + (({mcu[159:152], 8'b0} * 24'h08e)) + (({mcu[167:160], 8'b0} * 24'h08e)) + (({mcu[175:168], 8'b0} * 24'h08e)) + (({mcu[183:176], 8'b0} * 24'h08e)) + (({mcu[191:184], 8'b0} * 24'h08e)) + (({mcu[199:192], 8'b0} * 24'h031)) + (({mcu[207:200], 8'b0} * 24'h031)) + (({mcu[215:208], 8'b0} * 24'h031)) + (({mcu[223:216], 8'b0} * 24'h031)) + (({mcu[231:224], 8'b0} * 24'h031)) + (({mcu[239:232], 8'b0} * 24'h031)) + (({mcu[247:240], 8'b0} * 24'h031)) + (({mcu[255:248], 8'b0} * 24'h031)) + (({mcu[263:256], 8'b0} * -24'h031)) + (({mcu[271:264], 8'b0} * -24'h031)) + (({mcu[279:272], 8'b0} * -24'h031)) + (({mcu[287:280], 8'b0} * -24'h031)) + (({mcu[295:288], 8'b0} * -24'h031)) + (({mcu[303:296], 8'b0} * -24'h031)) + (({mcu[311:304], 8'b0} * -24'h031)) + (({mcu[319:312], 8'b0} * -24'h031)) + (({mcu[327:320], 8'b0} * -24'h08e)) + (({mcu[335:328], 8'b0} * -24'h08e)) + (({mcu[343:336], 8'b0} * -24'h08e)) + (({mcu[351:344], 8'b0} * -24'h08e)) + (({mcu[359:352], 8'b0} * -24'h08e)) + (({mcu[367:360], 8'b0} * -24'h08e)) + (({mcu[375:368], 8'b0} * -24'h08e)) + (({mcu[383:376], 8'b0} * -24'h08e)) + (({mcu[391:384], 8'b0} * -24'h0d4)) + (({mcu[399:392], 8'b0} * -24'h0d4)) + (({mcu[407:400], 8'b0} * -24'h0d4)) + (({mcu[415:408], 8'b0} * -24'h0d4)) + (({mcu[423:416], 8'b0} * -24'h0d4)) + (({mcu[431:424], 8'b0} * -24'h0d4)) + (({mcu[439:432], 8'b0} * -24'h0d4)) + (({mcu[447:440], 8'b0} * -24'h0d4)) + (({mcu[455:448], 8'b0} * -24'h0fb)) + (({mcu[463:456], 8'b0} * -24'h0fb)) + (({mcu[471:464], 8'b0} * -24'h0fb)) + (({mcu[479:472], 8'b0} * -24'h0fb)) + (({mcu[487:480], 8'b0} * -24'h0fb)) + (({mcu[495:488], 8'b0} * -24'h0fb)) + (({mcu[503:496], 8'b0} * -24'h0fb)) + (({mcu[511:504], 8'b0} * -24'h0fb));
	wire[47:0] cos11_term = (({mcu[7:0], 8'b0} * 24'h0f6)) + (({mcu[15:8], 8'b0} * 24'h0d0)) + (({mcu[23:16], 8'b0} * 24'h08b)) + (({mcu[31:24], 8'b0} * 24'h030)) + (({mcu[39:32], 8'b0} * -24'h030)) + (({mcu[47:40], 8'b0} * -24'h08b)) + (({mcu[55:48], 8'b0} * -24'h0d0)) + (({mcu[63:56], 8'b0} * -24'h0f6)) + (({mcu[71:64], 8'b0} * 24'h0d0)) + (({mcu[79:72], 8'b0} * 24'h0b0)) + (({mcu[87:80], 8'b0} * 24'h076)) + (({mcu[95:88], 8'b0} * 24'h029)) + (({mcu[103:96], 8'b0} * -24'h029)) + (({mcu[111:104], 8'b0} * -24'h076)) + (({mcu[119:112], 8'b0} * -24'h0b0)) + (({mcu[127:120], 8'b0} * -24'h0d0)) + (({mcu[135:128], 8'b0} * 24'h08b)) + (({mcu[143:136], 8'b0} * 24'h076)) + (({mcu[151:144], 8'b0} * 24'h04f)) + (({mcu[159:152], 8'b0} * 24'h01b)) + (({mcu[167:160], 8'b0} * -24'h01b)) + (({mcu[175:168], 8'b0} * -24'h04f)) + (({mcu[183:176], 8'b0} * -24'h076)) + (({mcu[191:184], 8'b0} * -24'h08b)) + (({mcu[199:192], 8'b0} * 24'h030)) + (({mcu[207:200], 8'b0} * 24'h029)) + (({mcu[215:208], 8'b0} * 24'h01b)) + (({mcu[223:216], 8'b0} * 24'h009)) + (({mcu[231:224], 8'b0} * -24'h009)) + (({mcu[239:232], 8'b0} * -24'h01b)) + (({mcu[247:240], 8'b0} * -24'h029)) + (({mcu[255:248], 8'b0} * -24'h030)) + (({mcu[263:256], 8'b0} * -24'h030)) + (({mcu[271:264], 8'b0} * -24'h029)) + (({mcu[279:272], 8'b0} * -24'h01b)) + (({mcu[287:280], 8'b0} * -24'h009)) + (({mcu[295:288], 8'b0} * 24'h009)) + (({mcu[303:296], 8'b0} * 24'h01b)) + (({mcu[311:304], 8'b0} * 24'h029)) + (({mcu[319:312], 8'b0} * 24'h030)) + (({mcu[327:320], 8'b0} * -24'h08b)) + (({mcu[335:328], 8'b0} * -24'h076)) + (({mcu[343:336], 8'b0} * -24'h04f)) + (({mcu[351:344], 8'b0} * -24'h01b)) + (({mcu[359:352], 8'b0} * 24'h01b)) + (({mcu[367:360], 8'b0} * 24'h04f)) + (({mcu[375:368], 8'b0} * 24'h076)) + (({mcu[383:376], 8'b0} * 24'h08b)) + (({mcu[391:384], 8'b0} * -24'h0d0)) + (({mcu[399:392], 8'b0} * -24'h0b0)) + (({mcu[407:400], 8'b0} * -24'h076)) + (({mcu[415:408], 8'b0} * -24'h029)) + (({mcu[423:416], 8'b0} * 24'h029)) + (({mcu[431:424], 8'b0} * 24'h076)) + (({mcu[439:432], 8'b0} * 24'h0b0)) + (({mcu[447:440], 8'b0} * 24'h0d0)) + (({mcu[455:448], 8'b0} * -24'h0f6)) + (({mcu[463:456], 8'b0} * -24'h0d0)) + (({mcu[471:464], 8'b0} * -24'h08b)) + (({mcu[479:472], 8'b0} * -24'h030)) + (({mcu[487:480], 8'b0} * 24'h030)) + (({mcu[495:488], 8'b0} * 24'h08b)) + (({mcu[503:496], 8'b0} * 24'h0d0)) + (({mcu[511:504], 8'b0} * 24'h0f6));
	wire[47:0] cos12_term = (({mcu[7:0], 8'b0} * 24'h0e7)) + (({mcu[15:8], 8'b0} * 24'h060)) + (({mcu[23:16], 8'b0} * -24'h060)) + (({mcu[31:24], 8'b0} * -24'h0e7)) + (({mcu[39:32], 8'b0} * -24'h0e7)) + (({mcu[47:40], 8'b0} * -24'h060)) + (({mcu[55:48], 8'b0} * 24'h060)) + (({mcu[63:56], 8'b0} * 24'h0e7)) + (({mcu[71:64], 8'b0} * 24'h0c4)) + (({mcu[79:72], 8'b0} * 24'h051)) + (({mcu[87:80], 8'b0} * -24'h051)) + (({mcu[95:88], 8'b0} * -24'h0c4)) + (({mcu[103:96], 8'b0} * -24'h0c4)) + (({mcu[111:104], 8'b0} * -24'h051)) + (({mcu[119:112], 8'b0} * 24'h051)) + (({mcu[127:120], 8'b0} * 24'h0c4)) + (({mcu[135:128], 8'b0} * 24'h083)) + (({mcu[143:136], 8'b0} * 24'h036)) + (({mcu[151:144], 8'b0} * -24'h036)) + (({mcu[159:152], 8'b0} * -24'h083)) + (({mcu[167:160], 8'b0} * -24'h083)) + (({mcu[175:168], 8'b0} * -24'h036)) + (({mcu[183:176], 8'b0} * 24'h036)) + (({mcu[191:184], 8'b0} * 24'h083)) + (({mcu[199:192], 8'b0} * 24'h02e)) + (({mcu[207:200], 8'b0} * 24'h013)) + (({mcu[215:208], 8'b0} * -24'h013)) + (({mcu[223:216], 8'b0} * -24'h02e)) + (({mcu[231:224], 8'b0} * -24'h02e)) + (({mcu[239:232], 8'b0} * -24'h013)) + (({mcu[247:240], 8'b0} * 24'h013)) + (({mcu[255:248], 8'b0} * 24'h02e)) + (({mcu[263:256], 8'b0} * -24'h02e)) + (({mcu[271:264], 8'b0} * -24'h013)) + (({mcu[279:272], 8'b0} * 24'h013)) + (({mcu[287:280], 8'b0} * 24'h02e)) + (({mcu[295:288], 8'b0} * 24'h02e)) + (({mcu[303:296], 8'b0} * 24'h013)) + (({mcu[311:304], 8'b0} * -24'h013)) + (({mcu[319:312], 8'b0} * -24'h02e)) + (({mcu[327:320], 8'b0} * -24'h083)) + (({mcu[335:328], 8'b0} * -24'h036)) + (({mcu[343:336], 8'b0} * 24'h036)) + (({mcu[351:344], 8'b0} * 24'h083)) + (({mcu[359:352], 8'b0} * 24'h083)) + (({mcu[367:360], 8'b0} * 24'h036)) + (({mcu[375:368], 8'b0} * -24'h036)) + (({mcu[383:376], 8'b0} * -24'h083)) + (({mcu[391:384], 8'b0} * -24'h0c4)) + (({mcu[399:392], 8'b0} * -24'h051)) + (({mcu[407:400], 8'b0} * 24'h051)) + (({mcu[415:408], 8'b0} * 24'h0c4)) + (({mcu[423:416], 8'b0} * 24'h0c4)) + (({mcu[431:424], 8'b0} * 24'h051)) + (({mcu[439:432], 8'b0} * -24'h051)) + (({mcu[447:440], 8'b0} * -24'h0c4)) + (({mcu[455:448], 8'b0} * -24'h0e7)) + (({mcu[463:456], 8'b0} * -24'h060)) + (({mcu[471:464], 8'b0} * 24'h060)) + (({mcu[479:472], 8'b0} * 24'h0e7)) + (({mcu[487:480], 8'b0} * 24'h0e7)) + (({mcu[495:488], 8'b0} * 24'h060)) + (({mcu[503:496], 8'b0} * -24'h060)) + (({mcu[511:504], 8'b0} * -24'h0e7));
	wire[47:0] cos13_term = (({mcu[7:0], 8'b0} * 24'h0d0)) + (({mcu[15:8], 8'b0} * -24'h030)) + (({mcu[23:16], 8'b0} * -24'h0f6)) + (({mcu[31:24], 8'b0} * -24'h08b)) + (({mcu[39:32], 8'b0} * 24'h08b)) + (({mcu[47:40], 8'b0} * 24'h0f6)) + (({mcu[55:48], 8'b0} * 24'h030)) + (({mcu[63:56], 8'b0} * -24'h0d0)) + (({mcu[71:64], 8'b0} * 24'h0b0)) + (({mcu[79:72], 8'b0} * -24'h029)) + (({mcu[87:80], 8'b0} * -24'h0d0)) + (({mcu[95:88], 8'b0} * -24'h076)) + (({mcu[103:96], 8'b0} * 24'h076)) + (({mcu[111:104], 8'b0} * 24'h0d0)) + (({mcu[119:112], 8'b0} * 24'h029)) + (({mcu[127:120], 8'b0} * -24'h0b0)) + (({mcu[135:128], 8'b0} * 24'h076)) + (({mcu[143:136], 8'b0} * -24'h01b)) + (({mcu[151:144], 8'b0} * -24'h08b)) + (({mcu[159:152], 8'b0} * -24'h04f)) + (({mcu[167:160], 8'b0} * 24'h04f)) + (({mcu[175:168], 8'b0} * 24'h08b)) + (({mcu[183:176], 8'b0} * 24'h01b)) + (({mcu[191:184], 8'b0} * -24'h076)) + (({mcu[199:192], 8'b0} * 24'h029)) + (({mcu[207:200], 8'b0} * -24'h009)) + (({mcu[215:208], 8'b0} * -24'h030)) + (({mcu[223:216], 8'b0} * -24'h01b)) + (({mcu[231:224], 8'b0} * 24'h01b)) + (({mcu[239:232], 8'b0} * 24'h030)) + (({mcu[247:240], 8'b0} * 24'h009)) + (({mcu[255:248], 8'b0} * -24'h029)) + (({mcu[263:256], 8'b0} * -24'h029)) + (({mcu[271:264], 8'b0} * 24'h009)) + (({mcu[279:272], 8'b0} * 24'h030)) + (({mcu[287:280], 8'b0} * 24'h01b)) + (({mcu[295:288], 8'b0} * -24'h01b)) + (({mcu[303:296], 8'b0} * -24'h030)) + (({mcu[311:304], 8'b0} * -24'h009)) + (({mcu[319:312], 8'b0} * 24'h029)) + (({mcu[327:320], 8'b0} * -24'h076)) + (({mcu[335:328], 8'b0} * 24'h01b)) + (({mcu[343:336], 8'b0} * 24'h08b)) + (({mcu[351:344], 8'b0} * 24'h04f)) + (({mcu[359:352], 8'b0} * -24'h04f)) + (({mcu[367:360], 8'b0} * -24'h08b)) + (({mcu[375:368], 8'b0} * -24'h01b)) + (({mcu[383:376], 8'b0} * 24'h076)) + (({mcu[391:384], 8'b0} * -24'h0b0)) + (({mcu[399:392], 8'b0} * 24'h029)) + (({mcu[407:400], 8'b0} * 24'h0d0)) + (({mcu[415:408], 8'b0} * 24'h076)) + (({mcu[423:416], 8'b0} * -24'h076)) + (({mcu[431:424], 8'b0} * -24'h0d0)) + (({mcu[439:432], 8'b0} * -24'h029)) + (({mcu[447:440], 8'b0} * 24'h0b0)) + (({mcu[455:448], 8'b0} * -24'h0d0)) + (({mcu[463:456], 8'b0} * 24'h030)) + (({mcu[471:464], 8'b0} * 24'h0f6)) + (({mcu[479:472], 8'b0} * 24'h08b)) + (({mcu[487:480], 8'b0} * -24'h08b)) + (({mcu[495:488], 8'b0} * -24'h0f6)) + (({mcu[503:496], 8'b0} * -24'h030)) + (({mcu[511:504], 8'b0} * 24'h0d0));
	wire[47:0] cos14_term = (({mcu[7:0], 8'b0} * 24'h0b1)) + (({mcu[15:8], 8'b0} * -24'h0b1)) + (({mcu[23:16], 8'b0} * -24'h0b1)) + (({mcu[31:24], 8'b0} * 24'h0b1)) + (({mcu[39:32], 8'b0} * 24'h0b1)) + (({mcu[47:40], 8'b0} * -24'h0b1)) + (({mcu[55:48], 8'b0} * -24'h0b1)) + (({mcu[63:56], 8'b0} * 24'h0b1)) + (({mcu[71:64], 8'b0} * 24'h096)) + (({mcu[79:72], 8'b0} * -24'h096)) + (({mcu[87:80], 8'b0} * -24'h096)) + (({mcu[95:88], 8'b0} * 24'h096)) + (({mcu[103:96], 8'b0} * 24'h096)) + (({mcu[111:104], 8'b0} * -24'h096)) + (({mcu[119:112], 8'b0} * -24'h096)) + (({mcu[127:120], 8'b0} * 24'h096)) + (({mcu[135:128], 8'b0} * 24'h064)) + (({mcu[143:136], 8'b0} * -24'h064)) + (({mcu[151:144], 8'b0} * -24'h064)) + (({mcu[159:152], 8'b0} * 24'h064)) + (({mcu[167:160], 8'b0} * 24'h064)) + (({mcu[175:168], 8'b0} * -24'h064)) + (({mcu[183:176], 8'b0} * -24'h064)) + (({mcu[191:184], 8'b0} * 24'h064)) + (({mcu[199:192], 8'b0} * 24'h023)) + (({mcu[207:200], 8'b0} * -24'h023)) + (({mcu[215:208], 8'b0} * -24'h023)) + (({mcu[223:216], 8'b0} * 24'h023)) + (({mcu[231:224], 8'b0} * 24'h023)) + (({mcu[239:232], 8'b0} * -24'h023)) + (({mcu[247:240], 8'b0} * -24'h023)) + (({mcu[255:248], 8'b0} * 24'h023)) + (({mcu[263:256], 8'b0} * -24'h023)) + (({mcu[271:264], 8'b0} * 24'h023)) + (({mcu[279:272], 8'b0} * 24'h023)) + (({mcu[287:280], 8'b0} * -24'h023)) + (({mcu[295:288], 8'b0} * -24'h023)) + (({mcu[303:296], 8'b0} * 24'h023)) + (({mcu[311:304], 8'b0} * 24'h023)) + (({mcu[319:312], 8'b0} * -24'h023)) + (({mcu[327:320], 8'b0} * -24'h064)) + (({mcu[335:328], 8'b0} * 24'h064)) + (({mcu[343:336], 8'b0} * 24'h064)) + (({mcu[351:344], 8'b0} * -24'h064)) + (({mcu[359:352], 8'b0} * -24'h064)) + (({mcu[367:360], 8'b0} * 24'h064)) + (({mcu[375:368], 8'b0} * 24'h064)) + (({mcu[383:376], 8'b0} * -24'h064)) + (({mcu[391:384], 8'b0} * -24'h096)) + (({mcu[399:392], 8'b0} * 24'h096)) + (({mcu[407:400], 8'b0} * 24'h096)) + (({mcu[415:408], 8'b0} * -24'h096)) + (({mcu[423:416], 8'b0} * -24'h096)) + (({mcu[431:424], 8'b0} * 24'h096)) + (({mcu[439:432], 8'b0} * 24'h096)) + (({mcu[447:440], 8'b0} * -24'h096)) + (({mcu[455:448], 8'b0} * -24'h0b1)) + (({mcu[463:456], 8'b0} * 24'h0b1)) + (({mcu[471:464], 8'b0} * 24'h0b1)) + (({mcu[479:472], 8'b0} * -24'h0b1)) + (({mcu[487:480], 8'b0} * -24'h0b1)) + (({mcu[495:488], 8'b0} * 24'h0b1)) + (({mcu[503:496], 8'b0} * 24'h0b1)) + (({mcu[511:504], 8'b0} * -24'h0b1));
	wire[47:0] cos15_term = (({mcu[7:0], 8'b0} * 24'h08b)) + (({mcu[15:8], 8'b0} * -24'h0f6)) + (({mcu[23:16], 8'b0} * 24'h030)) + (({mcu[31:24], 8'b0} * 24'h0d0)) + (({mcu[39:32], 8'b0} * -24'h0d0)) + (({mcu[47:40], 8'b0} * -24'h030)) + (({mcu[55:48], 8'b0} * 24'h0f6)) + (({mcu[63:56], 8'b0} * -24'h08b)) + (({mcu[71:64], 8'b0} * 24'h076)) + (({mcu[79:72], 8'b0} * -24'h0d0)) + (({mcu[87:80], 8'b0} * 24'h029)) + (({mcu[95:88], 8'b0} * 24'h0b0)) + (({mcu[103:96], 8'b0} * -24'h0b0)) + (({mcu[111:104], 8'b0} * -24'h029)) + (({mcu[119:112], 8'b0} * 24'h0d0)) + (({mcu[127:120], 8'b0} * -24'h076)) + (({mcu[135:128], 8'b0} * 24'h04f)) + (({mcu[143:136], 8'b0} * -24'h08b)) + (({mcu[151:144], 8'b0} * 24'h01b)) + (({mcu[159:152], 8'b0} * 24'h076)) + (({mcu[167:160], 8'b0} * -24'h076)) + (({mcu[175:168], 8'b0} * -24'h01b)) + (({mcu[183:176], 8'b0} * 24'h08b)) + (({mcu[191:184], 8'b0} * -24'h04f)) + (({mcu[199:192], 8'b0} * 24'h01b)) + (({mcu[207:200], 8'b0} * -24'h030)) + (({mcu[215:208], 8'b0} * 24'h009)) + (({mcu[223:216], 8'b0} * 24'h029)) + (({mcu[231:224], 8'b0} * -24'h029)) + (({mcu[239:232], 8'b0} * -24'h009)) + (({mcu[247:240], 8'b0} * 24'h030)) + (({mcu[255:248], 8'b0} * -24'h01b)) + (({mcu[263:256], 8'b0} * -24'h01b)) + (({mcu[271:264], 8'b0} * 24'h030)) + (({mcu[279:272], 8'b0} * -24'h009)) + (({mcu[287:280], 8'b0} * -24'h029)) + (({mcu[295:288], 8'b0} * 24'h029)) + (({mcu[303:296], 8'b0} * 24'h009)) + (({mcu[311:304], 8'b0} * -24'h030)) + (({mcu[319:312], 8'b0} * 24'h01b)) + (({mcu[327:320], 8'b0} * -24'h04f)) + (({mcu[335:328], 8'b0} * 24'h08b)) + (({mcu[343:336], 8'b0} * -24'h01b)) + (({mcu[351:344], 8'b0} * -24'h076)) + (({mcu[359:352], 8'b0} * 24'h076)) + (({mcu[367:360], 8'b0} * 24'h01b)) + (({mcu[375:368], 8'b0} * -24'h08b)) + (({mcu[383:376], 8'b0} * 24'h04f)) + (({mcu[391:384], 8'b0} * -24'h076)) + (({mcu[399:392], 8'b0} * 24'h0d0)) + (({mcu[407:400], 8'b0} * -24'h029)) + (({mcu[415:408], 8'b0} * -24'h0b0)) + (({mcu[423:416], 8'b0} * 24'h0b0)) + (({mcu[431:424], 8'b0} * 24'h029)) + (({mcu[439:432], 8'b0} * -24'h0d0)) + (({mcu[447:440], 8'b0} * 24'h076)) + (({mcu[455:448], 8'b0} * -24'h08b)) + (({mcu[463:456], 8'b0} * 24'h0f6)) + (({mcu[471:464], 8'b0} * -24'h030)) + (({mcu[479:472], 8'b0} * -24'h0d0)) + (({mcu[487:480], 8'b0} * 24'h0d0)) + (({mcu[495:488], 8'b0} * 24'h030)) + (({mcu[503:496], 8'b0} * -24'h0f6)) + (({mcu[511:504], 8'b0} * 24'h08b));
	wire[47:0] cos16_term = (({mcu[7:0], 8'b0} * 24'h060)) + (({mcu[15:8], 8'b0} * -24'h0e7)) + (({mcu[23:16], 8'b0} * 24'h0e7)) + (({mcu[31:24], 8'b0} * -24'h060)) + (({mcu[39:32], 8'b0} * -24'h060)) + (({mcu[47:40], 8'b0} * 24'h0e7)) + (({mcu[55:48], 8'b0} * -24'h0e7)) + (({mcu[63:56], 8'b0} * 24'h060)) + (({mcu[71:64], 8'b0} * 24'h051)) + (({mcu[79:72], 8'b0} * -24'h0c4)) + (({mcu[87:80], 8'b0} * 24'h0c4)) + (({mcu[95:88], 8'b0} * -24'h051)) + (({mcu[103:96], 8'b0} * -24'h051)) + (({mcu[111:104], 8'b0} * 24'h0c4)) + (({mcu[119:112], 8'b0} * -24'h0c4)) + (({mcu[127:120], 8'b0} * 24'h051)) + (({mcu[135:128], 8'b0} * 24'h036)) + (({mcu[143:136], 8'b0} * -24'h083)) + (({mcu[151:144], 8'b0} * 24'h083)) + (({mcu[159:152], 8'b0} * -24'h036)) + (({mcu[167:160], 8'b0} * -24'h036)) + (({mcu[175:168], 8'b0} * 24'h083)) + (({mcu[183:176], 8'b0} * -24'h083)) + (({mcu[191:184], 8'b0} * 24'h036)) + (({mcu[199:192], 8'b0} * 24'h013)) + (({mcu[207:200], 8'b0} * -24'h02e)) + (({mcu[215:208], 8'b0} * 24'h02e)) + (({mcu[223:216], 8'b0} * -24'h013)) + (({mcu[231:224], 8'b0} * -24'h013)) + (({mcu[239:232], 8'b0} * 24'h02e)) + (({mcu[247:240], 8'b0} * -24'h02e)) + (({mcu[255:248], 8'b0} * 24'h013)) + (({mcu[263:256], 8'b0} * -24'h013)) + (({mcu[271:264], 8'b0} * 24'h02e)) + (({mcu[279:272], 8'b0} * -24'h02e)) + (({mcu[287:280], 8'b0} * 24'h013)) + (({mcu[295:288], 8'b0} * 24'h013)) + (({mcu[303:296], 8'b0} * -24'h02e)) + (({mcu[311:304], 8'b0} * 24'h02e)) + (({mcu[319:312], 8'b0} * -24'h013)) + (({mcu[327:320], 8'b0} * -24'h036)) + (({mcu[335:328], 8'b0} * 24'h083)) + (({mcu[343:336], 8'b0} * -24'h083)) + (({mcu[351:344], 8'b0} * 24'h036)) + (({mcu[359:352], 8'b0} * 24'h036)) + (({mcu[367:360], 8'b0} * -24'h083)) + (({mcu[375:368], 8'b0} * 24'h083)) + (({mcu[383:376], 8'b0} * -24'h036)) + (({mcu[391:384], 8'b0} * -24'h051)) + (({mcu[399:392], 8'b0} * 24'h0c4)) + (({mcu[407:400], 8'b0} * -24'h0c4)) + (({mcu[415:408], 8'b0} * 24'h051)) + (({mcu[423:416], 8'b0} * 24'h051)) + (({mcu[431:424], 8'b0} * -24'h0c4)) + (({mcu[439:432], 8'b0} * 24'h0c4)) + (({mcu[447:440], 8'b0} * -24'h051)) + (({mcu[455:448], 8'b0} * -24'h060)) + (({mcu[463:456], 8'b0} * 24'h0e7)) + (({mcu[471:464], 8'b0} * -24'h0e7)) + (({mcu[479:472], 8'b0} * 24'h060)) + (({mcu[487:480], 8'b0} * 24'h060)) + (({mcu[495:488], 8'b0} * -24'h0e7)) + (({mcu[503:496], 8'b0} * 24'h0e7)) + (({mcu[511:504], 8'b0} * -24'h060));
	wire[47:0] cos17_term = (({mcu[7:0], 8'b0} * 24'h030)) + (({mcu[15:8], 8'b0} * -24'h08b)) + (({mcu[23:16], 8'b0} * 24'h0d0)) + (({mcu[31:24], 8'b0} * -24'h0f6)) + (({mcu[39:32], 8'b0} * 24'h0f6)) + (({mcu[47:40], 8'b0} * -24'h0d0)) + (({mcu[55:48], 8'b0} * 24'h08b)) + (({mcu[63:56], 8'b0} * -24'h030)) + (({mcu[71:64], 8'b0} * 24'h029)) + (({mcu[79:72], 8'b0} * -24'h076)) + (({mcu[87:80], 8'b0} * 24'h0b0)) + (({mcu[95:88], 8'b0} * -24'h0d0)) + (({mcu[103:96], 8'b0} * 24'h0d0)) + (({mcu[111:104], 8'b0} * -24'h0b0)) + (({mcu[119:112], 8'b0} * 24'h076)) + (({mcu[127:120], 8'b0} * -24'h029)) + (({mcu[135:128], 8'b0} * 24'h01b)) + (({mcu[143:136], 8'b0} * -24'h04f)) + (({mcu[151:144], 8'b0} * 24'h076)) + (({mcu[159:152], 8'b0} * -24'h08b)) + (({mcu[167:160], 8'b0} * 24'h08b)) + (({mcu[175:168], 8'b0} * -24'h076)) + (({mcu[183:176], 8'b0} * 24'h04f)) + (({mcu[191:184], 8'b0} * -24'h01b)) + (({mcu[199:192], 8'b0} * 24'h009)) + (({mcu[207:200], 8'b0} * -24'h01b)) + (({mcu[215:208], 8'b0} * 24'h029)) + (({mcu[223:216], 8'b0} * -24'h030)) + (({mcu[231:224], 8'b0} * 24'h030)) + (({mcu[239:232], 8'b0} * -24'h029)) + (({mcu[247:240], 8'b0} * 24'h01b)) + (({mcu[255:248], 8'b0} * -24'h009)) + (({mcu[263:256], 8'b0} * -24'h009)) + (({mcu[271:264], 8'b0} * 24'h01b)) + (({mcu[279:272], 8'b0} * -24'h029)) + (({mcu[287:280], 8'b0} * 24'h030)) + (({mcu[295:288], 8'b0} * -24'h030)) + (({mcu[303:296], 8'b0} * 24'h029)) + (({mcu[311:304], 8'b0} * -24'h01b)) + (({mcu[319:312], 8'b0} * 24'h009)) + (({mcu[327:320], 8'b0} * -24'h01b)) + (({mcu[335:328], 8'b0} * 24'h04f)) + (({mcu[343:336], 8'b0} * -24'h076)) + (({mcu[351:344], 8'b0} * 24'h08b)) + (({mcu[359:352], 8'b0} * -24'h08b)) + (({mcu[367:360], 8'b0} * 24'h076)) + (({mcu[375:368], 8'b0} * -24'h04f)) + (({mcu[383:376], 8'b0} * 24'h01b)) + (({mcu[391:384], 8'b0} * -24'h029)) + (({mcu[399:392], 8'b0} * 24'h076)) + (({mcu[407:400], 8'b0} * -24'h0b0)) + (({mcu[415:408], 8'b0} * 24'h0d0)) + (({mcu[423:416], 8'b0} * -24'h0d0)) + (({mcu[431:424], 8'b0} * 24'h0b0)) + (({mcu[439:432], 8'b0} * -24'h076)) + (({mcu[447:440], 8'b0} * 24'h029)) + (({mcu[455:448], 8'b0} * -24'h030)) + (({mcu[463:456], 8'b0} * 24'h08b)) + (({mcu[471:464], 8'b0} * -24'h0d0)) + (({mcu[479:472], 8'b0} * 24'h0f6)) + (({mcu[487:480], 8'b0} * -24'h0f6)) + (({mcu[495:488], 8'b0} * 24'h0d0)) + (({mcu[503:496], 8'b0} * -24'h08b)) + (({mcu[511:504], 8'b0} * 24'h030));
	wire[47:0] cos20_term = (({mcu[7:0], 8'b0} * 24'h0ec)) + (({mcu[15:8], 8'b0} * 24'h0ec)) + (({mcu[23:16], 8'b0} * 24'h0ec)) + (({mcu[31:24], 8'b0} * 24'h0ec)) + (({mcu[39:32], 8'b0} * 24'h0ec)) + (({mcu[47:40], 8'b0} * 24'h0ec)) + (({mcu[55:48], 8'b0} * 24'h0ec)) + (({mcu[63:56], 8'b0} * 24'h0ec)) + (({mcu[71:64], 8'b0} * 24'h062)) + (({mcu[79:72], 8'b0} * 24'h062)) + (({mcu[87:80], 8'b0} * 24'h062)) + (({mcu[95:88], 8'b0} * 24'h062)) + (({mcu[103:96], 8'b0} * 24'h062)) + (({mcu[111:104], 8'b0} * 24'h062)) + (({mcu[119:112], 8'b0} * 24'h062)) + (({mcu[127:120], 8'b0} * 24'h062)) + (({mcu[135:128], 8'b0} * -24'h062)) + (({mcu[143:136], 8'b0} * -24'h062)) + (({mcu[151:144], 8'b0} * -24'h062)) + (({mcu[159:152], 8'b0} * -24'h062)) + (({mcu[167:160], 8'b0} * -24'h062)) + (({mcu[175:168], 8'b0} * -24'h062)) + (({mcu[183:176], 8'b0} * -24'h062)) + (({mcu[191:184], 8'b0} * -24'h062)) + (({mcu[199:192], 8'b0} * -24'h0ec)) + (({mcu[207:200], 8'b0} * -24'h0ec)) + (({mcu[215:208], 8'b0} * -24'h0ec)) + (({mcu[223:216], 8'b0} * -24'h0ec)) + (({mcu[231:224], 8'b0} * -24'h0ec)) + (({mcu[239:232], 8'b0} * -24'h0ec)) + (({mcu[247:240], 8'b0} * -24'h0ec)) + (({mcu[255:248], 8'b0} * -24'h0ec)) + (({mcu[263:256], 8'b0} * -24'h0ec)) + (({mcu[271:264], 8'b0} * -24'h0ec)) + (({mcu[279:272], 8'b0} * -24'h0ec)) + (({mcu[287:280], 8'b0} * -24'h0ec)) + (({mcu[295:288], 8'b0} * -24'h0ec)) + (({mcu[303:296], 8'b0} * -24'h0ec)) + (({mcu[311:304], 8'b0} * -24'h0ec)) + (({mcu[319:312], 8'b0} * -24'h0ec)) + (({mcu[327:320], 8'b0} * -24'h062)) + (({mcu[335:328], 8'b0} * -24'h062)) + (({mcu[343:336], 8'b0} * -24'h062)) + (({mcu[351:344], 8'b0} * -24'h062)) + (({mcu[359:352], 8'b0} * -24'h062)) + (({mcu[367:360], 8'b0} * -24'h062)) + (({mcu[375:368], 8'b0} * -24'h062)) + (({mcu[383:376], 8'b0} * -24'h062)) + (({mcu[391:384], 8'b0} * 24'h062)) + (({mcu[399:392], 8'b0} * 24'h062)) + (({mcu[407:400], 8'b0} * 24'h062)) + (({mcu[415:408], 8'b0} * 24'h062)) + (({mcu[423:416], 8'b0} * 24'h062)) + (({mcu[431:424], 8'b0} * 24'h062)) + (({mcu[439:432], 8'b0} * 24'h062)) + (({mcu[447:440], 8'b0} * 24'h062)) + (({mcu[455:448], 8'b0} * 24'h0ec)) + (({mcu[463:456], 8'b0} * 24'h0ec)) + (({mcu[471:464], 8'b0} * 24'h0ec)) + (({mcu[479:472], 8'b0} * 24'h0ec)) + (({mcu[487:480], 8'b0} * 24'h0ec)) + (({mcu[495:488], 8'b0} * 24'h0ec)) + (({mcu[503:496], 8'b0} * 24'h0ec)) + (({mcu[511:504], 8'b0} * 24'h0ec));
	wire[47:0] cos21_term = (({mcu[7:0], 8'b0} * 24'h0e7)) + (({mcu[15:8], 8'b0} * 24'h0c4)) + (({mcu[23:16], 8'b0} * 24'h083)) + (({mcu[31:24], 8'b0} * 24'h02e)) + (({mcu[39:32], 8'b0} * -24'h02e)) + (({mcu[47:40], 8'b0} * -24'h083)) + (({mcu[55:48], 8'b0} * -24'h0c4)) + (({mcu[63:56], 8'b0} * -24'h0e7)) + (({mcu[71:64], 8'b0} * 24'h060)) + (({mcu[79:72], 8'b0} * 24'h051)) + (({mcu[87:80], 8'b0} * 24'h036)) + (({mcu[95:88], 8'b0} * 24'h013)) + (({mcu[103:96], 8'b0} * -24'h013)) + (({mcu[111:104], 8'b0} * -24'h036)) + (({mcu[119:112], 8'b0} * -24'h051)) + (({mcu[127:120], 8'b0} * -24'h060)) + (({mcu[135:128], 8'b0} * -24'h060)) + (({mcu[143:136], 8'b0} * -24'h051)) + (({mcu[151:144], 8'b0} * -24'h036)) + (({mcu[159:152], 8'b0} * -24'h013)) + (({mcu[167:160], 8'b0} * 24'h013)) + (({mcu[175:168], 8'b0} * 24'h036)) + (({mcu[183:176], 8'b0} * 24'h051)) + (({mcu[191:184], 8'b0} * 24'h060)) + (({mcu[199:192], 8'b0} * -24'h0e7)) + (({mcu[207:200], 8'b0} * -24'h0c4)) + (({mcu[215:208], 8'b0} * -24'h083)) + (({mcu[223:216], 8'b0} * -24'h02e)) + (({mcu[231:224], 8'b0} * 24'h02e)) + (({mcu[239:232], 8'b0} * 24'h083)) + (({mcu[247:240], 8'b0} * 24'h0c4)) + (({mcu[255:248], 8'b0} * 24'h0e7)) + (({mcu[263:256], 8'b0} * -24'h0e7)) + (({mcu[271:264], 8'b0} * -24'h0c4)) + (({mcu[279:272], 8'b0} * -24'h083)) + (({mcu[287:280], 8'b0} * -24'h02e)) + (({mcu[295:288], 8'b0} * 24'h02e)) + (({mcu[303:296], 8'b0} * 24'h083)) + (({mcu[311:304], 8'b0} * 24'h0c4)) + (({mcu[319:312], 8'b0} * 24'h0e7)) + (({mcu[327:320], 8'b0} * -24'h060)) + (({mcu[335:328], 8'b0} * -24'h051)) + (({mcu[343:336], 8'b0} * -24'h036)) + (({mcu[351:344], 8'b0} * -24'h013)) + (({mcu[359:352], 8'b0} * 24'h013)) + (({mcu[367:360], 8'b0} * 24'h036)) + (({mcu[375:368], 8'b0} * 24'h051)) + (({mcu[383:376], 8'b0} * 24'h060)) + (({mcu[391:384], 8'b0} * 24'h060)) + (({mcu[399:392], 8'b0} * 24'h051)) + (({mcu[407:400], 8'b0} * 24'h036)) + (({mcu[415:408], 8'b0} * 24'h013)) + (({mcu[423:416], 8'b0} * -24'h013)) + (({mcu[431:424], 8'b0} * -24'h036)) + (({mcu[439:432], 8'b0} * -24'h051)) + (({mcu[447:440], 8'b0} * -24'h060)) + (({mcu[455:448], 8'b0} * 24'h0e7)) + (({mcu[463:456], 8'b0} * 24'h0c4)) + (({mcu[471:464], 8'b0} * 24'h083)) + (({mcu[479:472], 8'b0} * 24'h02e)) + (({mcu[487:480], 8'b0} * -24'h02e)) + (({mcu[495:488], 8'b0} * -24'h083)) + (({mcu[503:496], 8'b0} * -24'h0c4)) + (({mcu[511:504], 8'b0} * -24'h0e7));
	wire[47:0] cos22_term = (({mcu[7:0], 8'b0} * 24'h0da)) + (({mcu[15:8], 8'b0} * 24'h05a)) + (({mcu[23:16], 8'b0} * -24'h05a)) + (({mcu[31:24], 8'b0} * -24'h0da)) + (({mcu[39:32], 8'b0} * -24'h0da)) + (({mcu[47:40], 8'b0} * -24'h05a)) + (({mcu[55:48], 8'b0} * 24'h05a)) + (({mcu[63:56], 8'b0} * 24'h0da)) + (({mcu[71:64], 8'b0} * 24'h05a)) + (({mcu[79:72], 8'b0} * 24'h025)) + (({mcu[87:80], 8'b0} * -24'h025)) + (({mcu[95:88], 8'b0} * -24'h05a)) + (({mcu[103:96], 8'b0} * -24'h05a)) + (({mcu[111:104], 8'b0} * -24'h025)) + (({mcu[119:112], 8'b0} * 24'h025)) + (({mcu[127:120], 8'b0} * 24'h05a)) + (({mcu[135:128], 8'b0} * -24'h05a)) + (({mcu[143:136], 8'b0} * -24'h025)) + (({mcu[151:144], 8'b0} * 24'h025)) + (({mcu[159:152], 8'b0} * 24'h05a)) + (({mcu[167:160], 8'b0} * 24'h05a)) + (({mcu[175:168], 8'b0} * 24'h025)) + (({mcu[183:176], 8'b0} * -24'h025)) + (({mcu[191:184], 8'b0} * -24'h05a)) + (({mcu[199:192], 8'b0} * -24'h0da)) + (({mcu[207:200], 8'b0} * -24'h05a)) + (({mcu[215:208], 8'b0} * 24'h05a)) + (({mcu[223:216], 8'b0} * 24'h0da)) + (({mcu[231:224], 8'b0} * 24'h0da)) + (({mcu[239:232], 8'b0} * 24'h05a)) + (({mcu[247:240], 8'b0} * -24'h05a)) + (({mcu[255:248], 8'b0} * -24'h0da)) + (({mcu[263:256], 8'b0} * -24'h0da)) + (({mcu[271:264], 8'b0} * -24'h05a)) + (({mcu[279:272], 8'b0} * 24'h05a)) + (({mcu[287:280], 8'b0} * 24'h0da)) + (({mcu[295:288], 8'b0} * 24'h0da)) + (({mcu[303:296], 8'b0} * 24'h05a)) + (({mcu[311:304], 8'b0} * -24'h05a)) + (({mcu[319:312], 8'b0} * -24'h0da)) + (({mcu[327:320], 8'b0} * -24'h05a)) + (({mcu[335:328], 8'b0} * -24'h025)) + (({mcu[343:336], 8'b0} * 24'h025)) + (({mcu[351:344], 8'b0} * 24'h05a)) + (({mcu[359:352], 8'b0} * 24'h05a)) + (({mcu[367:360], 8'b0} * 24'h025)) + (({mcu[375:368], 8'b0} * -24'h025)) + (({mcu[383:376], 8'b0} * -24'h05a)) + (({mcu[391:384], 8'b0} * 24'h05a)) + (({mcu[399:392], 8'b0} * 24'h025)) + (({mcu[407:400], 8'b0} * -24'h025)) + (({mcu[415:408], 8'b0} * -24'h05a)) + (({mcu[423:416], 8'b0} * -24'h05a)) + (({mcu[431:424], 8'b0} * -24'h025)) + (({mcu[439:432], 8'b0} * 24'h025)) + (({mcu[447:440], 8'b0} * 24'h05a)) + (({mcu[455:448], 8'b0} * 24'h0da)) + (({mcu[463:456], 8'b0} * 24'h05a)) + (({mcu[471:464], 8'b0} * -24'h05a)) + (({mcu[479:472], 8'b0} * -24'h0da)) + (({mcu[487:480], 8'b0} * -24'h0da)) + (({mcu[495:488], 8'b0} * -24'h05a)) + (({mcu[503:496], 8'b0} * 24'h05a)) + (({mcu[511:504], 8'b0} * 24'h0da));
	wire[47:0] cos23_term = (({mcu[7:0], 8'b0} * 24'h0c4)) + (({mcu[15:8], 8'b0} * -24'h02e)) + (({mcu[23:16], 8'b0} * -24'h0e7)) + (({mcu[31:24], 8'b0} * -24'h083)) + (({mcu[39:32], 8'b0} * 24'h083)) + (({mcu[47:40], 8'b0} * 24'h0e7)) + (({mcu[55:48], 8'b0} * 24'h02e)) + (({mcu[63:56], 8'b0} * -24'h0c4)) + (({mcu[71:64], 8'b0} * 24'h051)) + (({mcu[79:72], 8'b0} * -24'h013)) + (({mcu[87:80], 8'b0} * -24'h060)) + (({mcu[95:88], 8'b0} * -24'h036)) + (({mcu[103:96], 8'b0} * 24'h036)) + (({mcu[111:104], 8'b0} * 24'h060)) + (({mcu[119:112], 8'b0} * 24'h013)) + (({mcu[127:120], 8'b0} * -24'h051)) + (({mcu[135:128], 8'b0} * -24'h051)) + (({mcu[143:136], 8'b0} * 24'h013)) + (({mcu[151:144], 8'b0} * 24'h060)) + (({mcu[159:152], 8'b0} * 24'h036)) + (({mcu[167:160], 8'b0} * -24'h036)) + (({mcu[175:168], 8'b0} * -24'h060)) + (({mcu[183:176], 8'b0} * -24'h013)) + (({mcu[191:184], 8'b0} * 24'h051)) + (({mcu[199:192], 8'b0} * -24'h0c4)) + (({mcu[207:200], 8'b0} * 24'h02e)) + (({mcu[215:208], 8'b0} * 24'h0e7)) + (({mcu[223:216], 8'b0} * 24'h083)) + (({mcu[231:224], 8'b0} * -24'h083)) + (({mcu[239:232], 8'b0} * -24'h0e7)) + (({mcu[247:240], 8'b0} * -24'h02e)) + (({mcu[255:248], 8'b0} * 24'h0c4)) + (({mcu[263:256], 8'b0} * -24'h0c4)) + (({mcu[271:264], 8'b0} * 24'h02e)) + (({mcu[279:272], 8'b0} * 24'h0e7)) + (({mcu[287:280], 8'b0} * 24'h083)) + (({mcu[295:288], 8'b0} * -24'h083)) + (({mcu[303:296], 8'b0} * -24'h0e7)) + (({mcu[311:304], 8'b0} * -24'h02e)) + (({mcu[319:312], 8'b0} * 24'h0c4)) + (({mcu[327:320], 8'b0} * -24'h051)) + (({mcu[335:328], 8'b0} * 24'h013)) + (({mcu[343:336], 8'b0} * 24'h060)) + (({mcu[351:344], 8'b0} * 24'h036)) + (({mcu[359:352], 8'b0} * -24'h036)) + (({mcu[367:360], 8'b0} * -24'h060)) + (({mcu[375:368], 8'b0} * -24'h013)) + (({mcu[383:376], 8'b0} * 24'h051)) + (({mcu[391:384], 8'b0} * 24'h051)) + (({mcu[399:392], 8'b0} * -24'h013)) + (({mcu[407:400], 8'b0} * -24'h060)) + (({mcu[415:408], 8'b0} * -24'h036)) + (({mcu[423:416], 8'b0} * 24'h036)) + (({mcu[431:424], 8'b0} * 24'h060)) + (({mcu[439:432], 8'b0} * 24'h013)) + (({mcu[447:440], 8'b0} * -24'h051)) + (({mcu[455:448], 8'b0} * 24'h0c4)) + (({mcu[463:456], 8'b0} * -24'h02e)) + (({mcu[471:464], 8'b0} * -24'h0e7)) + (({mcu[479:472], 8'b0} * -24'h083)) + (({mcu[487:480], 8'b0} * 24'h083)) + (({mcu[495:488], 8'b0} * 24'h0e7)) + (({mcu[503:496], 8'b0} * 24'h02e)) + (({mcu[511:504], 8'b0} * -24'h0c4));
	wire[47:0] cos24_term = (({mcu[7:0], 8'b0} * 24'h0a7)) + (({mcu[15:8], 8'b0} * -24'h0a7)) + (({mcu[23:16], 8'b0} * -24'h0a7)) + (({mcu[31:24], 8'b0} * 24'h0a7)) + (({mcu[39:32], 8'b0} * 24'h0a7)) + (({mcu[47:40], 8'b0} * -24'h0a7)) + (({mcu[55:48], 8'b0} * -24'h0a7)) + (({mcu[63:56], 8'b0} * 24'h0a7)) + (({mcu[71:64], 8'b0} * 24'h045)) + (({mcu[79:72], 8'b0} * -24'h045)) + (({mcu[87:80], 8'b0} * -24'h045)) + (({mcu[95:88], 8'b0} * 24'h045)) + (({mcu[103:96], 8'b0} * 24'h045)) + (({mcu[111:104], 8'b0} * -24'h045)) + (({mcu[119:112], 8'b0} * -24'h045)) + (({mcu[127:120], 8'b0} * 24'h045)) + (({mcu[135:128], 8'b0} * -24'h045)) + (({mcu[143:136], 8'b0} * 24'h045)) + (({mcu[151:144], 8'b0} * 24'h045)) + (({mcu[159:152], 8'b0} * -24'h045)) + (({mcu[167:160], 8'b0} * -24'h045)) + (({mcu[175:168], 8'b0} * 24'h045)) + (({mcu[183:176], 8'b0} * 24'h045)) + (({mcu[191:184], 8'b0} * -24'h045)) + (({mcu[199:192], 8'b0} * -24'h0a7)) + (({mcu[207:200], 8'b0} * 24'h0a7)) + (({mcu[215:208], 8'b0} * 24'h0a7)) + (({mcu[223:216], 8'b0} * -24'h0a7)) + (({mcu[231:224], 8'b0} * -24'h0a7)) + (({mcu[239:232], 8'b0} * 24'h0a7)) + (({mcu[247:240], 8'b0} * 24'h0a7)) + (({mcu[255:248], 8'b0} * -24'h0a7)) + (({mcu[263:256], 8'b0} * -24'h0a7)) + (({mcu[271:264], 8'b0} * 24'h0a7)) + (({mcu[279:272], 8'b0} * 24'h0a7)) + (({mcu[287:280], 8'b0} * -24'h0a7)) + (({mcu[295:288], 8'b0} * -24'h0a7)) + (({mcu[303:296], 8'b0} * 24'h0a7)) + (({mcu[311:304], 8'b0} * 24'h0a7)) + (({mcu[319:312], 8'b0} * -24'h0a7)) + (({mcu[327:320], 8'b0} * -24'h045)) + (({mcu[335:328], 8'b0} * 24'h045)) + (({mcu[343:336], 8'b0} * 24'h045)) + (({mcu[351:344], 8'b0} * -24'h045)) + (({mcu[359:352], 8'b0} * -24'h045)) + (({mcu[367:360], 8'b0} * 24'h045)) + (({mcu[375:368], 8'b0} * 24'h045)) + (({mcu[383:376], 8'b0} * -24'h045)) + (({mcu[391:384], 8'b0} * 24'h045)) + (({mcu[399:392], 8'b0} * -24'h045)) + (({mcu[407:400], 8'b0} * -24'h045)) + (({mcu[415:408], 8'b0} * 24'h045)) + (({mcu[423:416], 8'b0} * 24'h045)) + (({mcu[431:424], 8'b0} * -24'h045)) + (({mcu[439:432], 8'b0} * -24'h045)) + (({mcu[447:440], 8'b0} * 24'h045)) + (({mcu[455:448], 8'b0} * 24'h0a7)) + (({mcu[463:456], 8'b0} * -24'h0a7)) + (({mcu[471:464], 8'b0} * -24'h0a7)) + (({mcu[479:472], 8'b0} * 24'h0a7)) + (({mcu[487:480], 8'b0} * 24'h0a7)) + (({mcu[495:488], 8'b0} * -24'h0a7)) + (({mcu[503:496], 8'b0} * -24'h0a7)) + (({mcu[511:504], 8'b0} * 24'h0a7));
	wire[47:0] cos25_term = (({mcu[7:0], 8'b0} * 24'h083)) + (({mcu[15:8], 8'b0} * -24'h0e7)) + (({mcu[23:16], 8'b0} * 24'h02e)) + (({mcu[31:24], 8'b0} * 24'h0c4)) + (({mcu[39:32], 8'b0} * -24'h0c4)) + (({mcu[47:40], 8'b0} * -24'h02e)) + (({mcu[55:48], 8'b0} * 24'h0e7)) + (({mcu[63:56], 8'b0} * -24'h083)) + (({mcu[71:64], 8'b0} * 24'h036)) + (({mcu[79:72], 8'b0} * -24'h060)) + (({mcu[87:80], 8'b0} * 24'h013)) + (({mcu[95:88], 8'b0} * 24'h051)) + (({mcu[103:96], 8'b0} * -24'h051)) + (({mcu[111:104], 8'b0} * -24'h013)) + (({mcu[119:112], 8'b0} * 24'h060)) + (({mcu[127:120], 8'b0} * -24'h036)) + (({mcu[135:128], 8'b0} * -24'h036)) + (({mcu[143:136], 8'b0} * 24'h060)) + (({mcu[151:144], 8'b0} * -24'h013)) + (({mcu[159:152], 8'b0} * -24'h051)) + (({mcu[167:160], 8'b0} * 24'h051)) + (({mcu[175:168], 8'b0} * 24'h013)) + (({mcu[183:176], 8'b0} * -24'h060)) + (({mcu[191:184], 8'b0} * 24'h036)) + (({mcu[199:192], 8'b0} * -24'h083)) + (({mcu[207:200], 8'b0} * 24'h0e7)) + (({mcu[215:208], 8'b0} * -24'h02e)) + (({mcu[223:216], 8'b0} * -24'h0c4)) + (({mcu[231:224], 8'b0} * 24'h0c4)) + (({mcu[239:232], 8'b0} * 24'h02e)) + (({mcu[247:240], 8'b0} * -24'h0e7)) + (({mcu[255:248], 8'b0} * 24'h083)) + (({mcu[263:256], 8'b0} * -24'h083)) + (({mcu[271:264], 8'b0} * 24'h0e7)) + (({mcu[279:272], 8'b0} * -24'h02e)) + (({mcu[287:280], 8'b0} * -24'h0c4)) + (({mcu[295:288], 8'b0} * 24'h0c4)) + (({mcu[303:296], 8'b0} * 24'h02e)) + (({mcu[311:304], 8'b0} * -24'h0e7)) + (({mcu[319:312], 8'b0} * 24'h083)) + (({mcu[327:320], 8'b0} * -24'h036)) + (({mcu[335:328], 8'b0} * 24'h060)) + (({mcu[343:336], 8'b0} * -24'h013)) + (({mcu[351:344], 8'b0} * -24'h051)) + (({mcu[359:352], 8'b0} * 24'h051)) + (({mcu[367:360], 8'b0} * 24'h013)) + (({mcu[375:368], 8'b0} * -24'h060)) + (({mcu[383:376], 8'b0} * 24'h036)) + (({mcu[391:384], 8'b0} * 24'h036)) + (({mcu[399:392], 8'b0} * -24'h060)) + (({mcu[407:400], 8'b0} * 24'h013)) + (({mcu[415:408], 8'b0} * 24'h051)) + (({mcu[423:416], 8'b0} * -24'h051)) + (({mcu[431:424], 8'b0} * -24'h013)) + (({mcu[439:432], 8'b0} * 24'h060)) + (({mcu[447:440], 8'b0} * -24'h036)) + (({mcu[455:448], 8'b0} * 24'h083)) + (({mcu[463:456], 8'b0} * -24'h0e7)) + (({mcu[471:464], 8'b0} * 24'h02e)) + (({mcu[479:472], 8'b0} * 24'h0c4)) + (({mcu[487:480], 8'b0} * -24'h0c4)) + (({mcu[495:488], 8'b0} * -24'h02e)) + (({mcu[503:496], 8'b0} * 24'h0e7)) + (({mcu[511:504], 8'b0} * -24'h083));
	wire[47:0] cos26_term = (({mcu[7:0], 8'b0} * 24'h05a)) + (({mcu[15:8], 8'b0} * -24'h0da)) + (({mcu[23:16], 8'b0} * 24'h0da)) + (({mcu[31:24], 8'b0} * -24'h05a)) + (({mcu[39:32], 8'b0} * -24'h05a)) + (({mcu[47:40], 8'b0} * 24'h0da)) + (({mcu[55:48], 8'b0} * -24'h0da)) + (({mcu[63:56], 8'b0} * 24'h05a)) + (({mcu[71:64], 8'b0} * 24'h025)) + (({mcu[79:72], 8'b0} * -24'h05a)) + (({mcu[87:80], 8'b0} * 24'h05a)) + (({mcu[95:88], 8'b0} * -24'h025)) + (({mcu[103:96], 8'b0} * -24'h025)) + (({mcu[111:104], 8'b0} * 24'h05a)) + (({mcu[119:112], 8'b0} * -24'h05a)) + (({mcu[127:120], 8'b0} * 24'h025)) + (({mcu[135:128], 8'b0} * -24'h025)) + (({mcu[143:136], 8'b0} * 24'h05a)) + (({mcu[151:144], 8'b0} * -24'h05a)) + (({mcu[159:152], 8'b0} * 24'h025)) + (({mcu[167:160], 8'b0} * 24'h025)) + (({mcu[175:168], 8'b0} * -24'h05a)) + (({mcu[183:176], 8'b0} * 24'h05a)) + (({mcu[191:184], 8'b0} * -24'h025)) + (({mcu[199:192], 8'b0} * -24'h05a)) + (({mcu[207:200], 8'b0} * 24'h0da)) + (({mcu[215:208], 8'b0} * -24'h0da)) + (({mcu[223:216], 8'b0} * 24'h05a)) + (({mcu[231:224], 8'b0} * 24'h05a)) + (({mcu[239:232], 8'b0} * -24'h0da)) + (({mcu[247:240], 8'b0} * 24'h0da)) + (({mcu[255:248], 8'b0} * -24'h05a)) + (({mcu[263:256], 8'b0} * -24'h05a)) + (({mcu[271:264], 8'b0} * 24'h0da)) + (({mcu[279:272], 8'b0} * -24'h0da)) + (({mcu[287:280], 8'b0} * 24'h05a)) + (({mcu[295:288], 8'b0} * 24'h05a)) + (({mcu[303:296], 8'b0} * -24'h0da)) + (({mcu[311:304], 8'b0} * 24'h0da)) + (({mcu[319:312], 8'b0} * -24'h05a)) + (({mcu[327:320], 8'b0} * -24'h025)) + (({mcu[335:328], 8'b0} * 24'h05a)) + (({mcu[343:336], 8'b0} * -24'h05a)) + (({mcu[351:344], 8'b0} * 24'h025)) + (({mcu[359:352], 8'b0} * 24'h025)) + (({mcu[367:360], 8'b0} * -24'h05a)) + (({mcu[375:368], 8'b0} * 24'h05a)) + (({mcu[383:376], 8'b0} * -24'h025)) + (({mcu[391:384], 8'b0} * 24'h025)) + (({mcu[399:392], 8'b0} * -24'h05a)) + (({mcu[407:400], 8'b0} * 24'h05a)) + (({mcu[415:408], 8'b0} * -24'h025)) + (({mcu[423:416], 8'b0} * -24'h025)) + (({mcu[431:424], 8'b0} * 24'h05a)) + (({mcu[439:432], 8'b0} * -24'h05a)) + (({mcu[447:440], 8'b0} * 24'h025)) + (({mcu[455:448], 8'b0} * 24'h05a)) + (({mcu[463:456], 8'b0} * -24'h0da)) + (({mcu[471:464], 8'b0} * 24'h0da)) + (({mcu[479:472], 8'b0} * -24'h05a)) + (({mcu[487:480], 8'b0} * -24'h05a)) + (({mcu[495:488], 8'b0} * 24'h0da)) + (({mcu[503:496], 8'b0} * -24'h0da)) + (({mcu[511:504], 8'b0} * 24'h05a));
	wire[47:0] cos27_term = (({mcu[7:0], 8'b0} * 24'h02e)) + (({mcu[15:8], 8'b0} * -24'h083)) + (({mcu[23:16], 8'b0} * 24'h0c4)) + (({mcu[31:24], 8'b0} * -24'h0e7)) + (({mcu[39:32], 8'b0} * 24'h0e7)) + (({mcu[47:40], 8'b0} * -24'h0c4)) + (({mcu[55:48], 8'b0} * 24'h083)) + (({mcu[63:56], 8'b0} * -24'h02e)) + (({mcu[71:64], 8'b0} * 24'h013)) + (({mcu[79:72], 8'b0} * -24'h036)) + (({mcu[87:80], 8'b0} * 24'h051)) + (({mcu[95:88], 8'b0} * -24'h060)) + (({mcu[103:96], 8'b0} * 24'h060)) + (({mcu[111:104], 8'b0} * -24'h051)) + (({mcu[119:112], 8'b0} * 24'h036)) + (({mcu[127:120], 8'b0} * -24'h013)) + (({mcu[135:128], 8'b0} * -24'h013)) + (({mcu[143:136], 8'b0} * 24'h036)) + (({mcu[151:144], 8'b0} * -24'h051)) + (({mcu[159:152], 8'b0} * 24'h060)) + (({mcu[167:160], 8'b0} * -24'h060)) + (({mcu[175:168], 8'b0} * 24'h051)) + (({mcu[183:176], 8'b0} * -24'h036)) + (({mcu[191:184], 8'b0} * 24'h013)) + (({mcu[199:192], 8'b0} * -24'h02e)) + (({mcu[207:200], 8'b0} * 24'h083)) + (({mcu[215:208], 8'b0} * -24'h0c4)) + (({mcu[223:216], 8'b0} * 24'h0e7)) + (({mcu[231:224], 8'b0} * -24'h0e7)) + (({mcu[239:232], 8'b0} * 24'h0c4)) + (({mcu[247:240], 8'b0} * -24'h083)) + (({mcu[255:248], 8'b0} * 24'h02e)) + (({mcu[263:256], 8'b0} * -24'h02e)) + (({mcu[271:264], 8'b0} * 24'h083)) + (({mcu[279:272], 8'b0} * -24'h0c4)) + (({mcu[287:280], 8'b0} * 24'h0e7)) + (({mcu[295:288], 8'b0} * -24'h0e7)) + (({mcu[303:296], 8'b0} * 24'h0c4)) + (({mcu[311:304], 8'b0} * -24'h083)) + (({mcu[319:312], 8'b0} * 24'h02e)) + (({mcu[327:320], 8'b0} * -24'h013)) + (({mcu[335:328], 8'b0} * 24'h036)) + (({mcu[343:336], 8'b0} * -24'h051)) + (({mcu[351:344], 8'b0} * 24'h060)) + (({mcu[359:352], 8'b0} * -24'h060)) + (({mcu[367:360], 8'b0} * 24'h051)) + (({mcu[375:368], 8'b0} * -24'h036)) + (({mcu[383:376], 8'b0} * 24'h013)) + (({mcu[391:384], 8'b0} * 24'h013)) + (({mcu[399:392], 8'b0} * -24'h036)) + (({mcu[407:400], 8'b0} * 24'h051)) + (({mcu[415:408], 8'b0} * -24'h060)) + (({mcu[423:416], 8'b0} * 24'h060)) + (({mcu[431:424], 8'b0} * -24'h051)) + (({mcu[439:432], 8'b0} * 24'h036)) + (({mcu[447:440], 8'b0} * -24'h013)) + (({mcu[455:448], 8'b0} * 24'h02e)) + (({mcu[463:456], 8'b0} * -24'h083)) + (({mcu[471:464], 8'b0} * 24'h0c4)) + (({mcu[479:472], 8'b0} * -24'h0e7)) + (({mcu[487:480], 8'b0} * 24'h0e7)) + (({mcu[495:488], 8'b0} * -24'h0c4)) + (({mcu[503:496], 8'b0} * 24'h083)) + (({mcu[511:504], 8'b0} * -24'h02e));
	wire[47:0] cos30_term = (({mcu[7:0], 8'b0} * 24'h0d4)) + (({mcu[15:8], 8'b0} * 24'h0d4)) + (({mcu[23:16], 8'b0} * 24'h0d4)) + (({mcu[31:24], 8'b0} * 24'h0d4)) + (({mcu[39:32], 8'b0} * 24'h0d4)) + (({mcu[47:40], 8'b0} * 24'h0d4)) + (({mcu[55:48], 8'b0} * 24'h0d4)) + (({mcu[63:56], 8'b0} * 24'h0d4)) + (({mcu[71:64], 8'b0} * -24'h031)) + (({mcu[79:72], 8'b0} * -24'h031)) + (({mcu[87:80], 8'b0} * -24'h031)) + (({mcu[95:88], 8'b0} * -24'h031)) + (({mcu[103:96], 8'b0} * -24'h031)) + (({mcu[111:104], 8'b0} * -24'h031)) + (({mcu[119:112], 8'b0} * -24'h031)) + (({mcu[127:120], 8'b0} * -24'h031)) + (({mcu[135:128], 8'b0} * -24'h0fb)) + (({mcu[143:136], 8'b0} * -24'h0fb)) + (({mcu[151:144], 8'b0} * -24'h0fb)) + (({mcu[159:152], 8'b0} * -24'h0fb)) + (({mcu[167:160], 8'b0} * -24'h0fb)) + (({mcu[175:168], 8'b0} * -24'h0fb)) + (({mcu[183:176], 8'b0} * -24'h0fb)) + (({mcu[191:184], 8'b0} * -24'h0fb)) + (({mcu[199:192], 8'b0} * -24'h08e)) + (({mcu[207:200], 8'b0} * -24'h08e)) + (({mcu[215:208], 8'b0} * -24'h08e)) + (({mcu[223:216], 8'b0} * -24'h08e)) + (({mcu[231:224], 8'b0} * -24'h08e)) + (({mcu[239:232], 8'b0} * -24'h08e)) + (({mcu[247:240], 8'b0} * -24'h08e)) + (({mcu[255:248], 8'b0} * -24'h08e)) + (({mcu[263:256], 8'b0} * 24'h08e)) + (({mcu[271:264], 8'b0} * 24'h08e)) + (({mcu[279:272], 8'b0} * 24'h08e)) + (({mcu[287:280], 8'b0} * 24'h08e)) + (({mcu[295:288], 8'b0} * 24'h08e)) + (({mcu[303:296], 8'b0} * 24'h08e)) + (({mcu[311:304], 8'b0} * 24'h08e)) + (({mcu[319:312], 8'b0} * 24'h08e)) + (({mcu[327:320], 8'b0} * 24'h0fb)) + (({mcu[335:328], 8'b0} * 24'h0fb)) + (({mcu[343:336], 8'b0} * 24'h0fb)) + (({mcu[351:344], 8'b0} * 24'h0fb)) + (({mcu[359:352], 8'b0} * 24'h0fb)) + (({mcu[367:360], 8'b0} * 24'h0fb)) + (({mcu[375:368], 8'b0} * 24'h0fb)) + (({mcu[383:376], 8'b0} * 24'h0fb)) + (({mcu[391:384], 8'b0} * 24'h031)) + (({mcu[399:392], 8'b0} * 24'h031)) + (({mcu[407:400], 8'b0} * 24'h031)) + (({mcu[415:408], 8'b0} * 24'h031)) + (({mcu[423:416], 8'b0} * 24'h031)) + (({mcu[431:424], 8'b0} * 24'h031)) + (({mcu[439:432], 8'b0} * 24'h031)) + (({mcu[447:440], 8'b0} * 24'h031)) + (({mcu[455:448], 8'b0} * -24'h0d4)) + (({mcu[463:456], 8'b0} * -24'h0d4)) + (({mcu[471:464], 8'b0} * -24'h0d4)) + (({mcu[479:472], 8'b0} * -24'h0d4)) + (({mcu[487:480], 8'b0} * -24'h0d4)) + (({mcu[495:488], 8'b0} * -24'h0d4)) + (({mcu[503:496], 8'b0} * -24'h0d4)) + (({mcu[511:504], 8'b0} * -24'h0d4));
	wire[47:0] cos31_term = (({mcu[7:0], 8'b0} * 24'h0d0)) + (({mcu[15:8], 8'b0} * 24'h0b0)) + (({mcu[23:16], 8'b0} * 24'h076)) + (({mcu[31:24], 8'b0} * 24'h029)) + (({mcu[39:32], 8'b0} * -24'h029)) + (({mcu[47:40], 8'b0} * -24'h076)) + (({mcu[55:48], 8'b0} * -24'h0b0)) + (({mcu[63:56], 8'b0} * -24'h0d0)) + (({mcu[71:64], 8'b0} * -24'h030)) + (({mcu[79:72], 8'b0} * -24'h029)) + (({mcu[87:80], 8'b0} * -24'h01b)) + (({mcu[95:88], 8'b0} * -24'h009)) + (({mcu[103:96], 8'b0} * 24'h009)) + (({mcu[111:104], 8'b0} * 24'h01b)) + (({mcu[119:112], 8'b0} * 24'h029)) + (({mcu[127:120], 8'b0} * 24'h030)) + (({mcu[135:128], 8'b0} * -24'h0f6)) + (({mcu[143:136], 8'b0} * -24'h0d0)) + (({mcu[151:144], 8'b0} * -24'h08b)) + (({mcu[159:152], 8'b0} * -24'h030)) + (({mcu[167:160], 8'b0} * 24'h030)) + (({mcu[175:168], 8'b0} * 24'h08b)) + (({mcu[183:176], 8'b0} * 24'h0d0)) + (({mcu[191:184], 8'b0} * 24'h0f6)) + (({mcu[199:192], 8'b0} * -24'h08b)) + (({mcu[207:200], 8'b0} * -24'h076)) + (({mcu[215:208], 8'b0} * -24'h04f)) + (({mcu[223:216], 8'b0} * -24'h01b)) + (({mcu[231:224], 8'b0} * 24'h01b)) + (({mcu[239:232], 8'b0} * 24'h04f)) + (({mcu[247:240], 8'b0} * 24'h076)) + (({mcu[255:248], 8'b0} * 24'h08b)) + (({mcu[263:256], 8'b0} * 24'h08b)) + (({mcu[271:264], 8'b0} * 24'h076)) + (({mcu[279:272], 8'b0} * 24'h04f)) + (({mcu[287:280], 8'b0} * 24'h01b)) + (({mcu[295:288], 8'b0} * -24'h01b)) + (({mcu[303:296], 8'b0} * -24'h04f)) + (({mcu[311:304], 8'b0} * -24'h076)) + (({mcu[319:312], 8'b0} * -24'h08b)) + (({mcu[327:320], 8'b0} * 24'h0f6)) + (({mcu[335:328], 8'b0} * 24'h0d0)) + (({mcu[343:336], 8'b0} * 24'h08b)) + (({mcu[351:344], 8'b0} * 24'h030)) + (({mcu[359:352], 8'b0} * -24'h030)) + (({mcu[367:360], 8'b0} * -24'h08b)) + (({mcu[375:368], 8'b0} * -24'h0d0)) + (({mcu[383:376], 8'b0} * -24'h0f6)) + (({mcu[391:384], 8'b0} * 24'h030)) + (({mcu[399:392], 8'b0} * 24'h029)) + (({mcu[407:400], 8'b0} * 24'h01b)) + (({mcu[415:408], 8'b0} * 24'h009)) + (({mcu[423:416], 8'b0} * -24'h009)) + (({mcu[431:424], 8'b0} * -24'h01b)) + (({mcu[439:432], 8'b0} * -24'h029)) + (({mcu[447:440], 8'b0} * -24'h030)) + (({mcu[455:448], 8'b0} * -24'h0d0)) + (({mcu[463:456], 8'b0} * -24'h0b0)) + (({mcu[471:464], 8'b0} * -24'h076)) + (({mcu[479:472], 8'b0} * -24'h029)) + (({mcu[487:480], 8'b0} * 24'h029)) + (({mcu[495:488], 8'b0} * 24'h076)) + (({mcu[503:496], 8'b0} * 24'h0b0)) + (({mcu[511:504], 8'b0} * 24'h0d0));
	wire[47:0] cos32_term = (({mcu[7:0], 8'b0} * 24'h0c4)) + (({mcu[15:8], 8'b0} * 24'h051)) + (({mcu[23:16], 8'b0} * -24'h051)) + (({mcu[31:24], 8'b0} * -24'h0c4)) + (({mcu[39:32], 8'b0} * -24'h0c4)) + (({mcu[47:40], 8'b0} * -24'h051)) + (({mcu[55:48], 8'b0} * 24'h051)) + (({mcu[63:56], 8'b0} * 24'h0c4)) + (({mcu[71:64], 8'b0} * -24'h02e)) + (({mcu[79:72], 8'b0} * -24'h013)) + (({mcu[87:80], 8'b0} * 24'h013)) + (({mcu[95:88], 8'b0} * 24'h02e)) + (({mcu[103:96], 8'b0} * 24'h02e)) + (({mcu[111:104], 8'b0} * 24'h013)) + (({mcu[119:112], 8'b0} * -24'h013)) + (({mcu[127:120], 8'b0} * -24'h02e)) + (({mcu[135:128], 8'b0} * -24'h0e7)) + (({mcu[143:136], 8'b0} * -24'h060)) + (({mcu[151:144], 8'b0} * 24'h060)) + (({mcu[159:152], 8'b0} * 24'h0e7)) + (({mcu[167:160], 8'b0} * 24'h0e7)) + (({mcu[175:168], 8'b0} * 24'h060)) + (({mcu[183:176], 8'b0} * -24'h060)) + (({mcu[191:184], 8'b0} * -24'h0e7)) + (({mcu[199:192], 8'b0} * -24'h083)) + (({mcu[207:200], 8'b0} * -24'h036)) + (({mcu[215:208], 8'b0} * 24'h036)) + (({mcu[223:216], 8'b0} * 24'h083)) + (({mcu[231:224], 8'b0} * 24'h083)) + (({mcu[239:232], 8'b0} * 24'h036)) + (({mcu[247:240], 8'b0} * -24'h036)) + (({mcu[255:248], 8'b0} * -24'h083)) + (({mcu[263:256], 8'b0} * 24'h083)) + (({mcu[271:264], 8'b0} * 24'h036)) + (({mcu[279:272], 8'b0} * -24'h036)) + (({mcu[287:280], 8'b0} * -24'h083)) + (({mcu[295:288], 8'b0} * -24'h083)) + (({mcu[303:296], 8'b0} * -24'h036)) + (({mcu[311:304], 8'b0} * 24'h036)) + (({mcu[319:312], 8'b0} * 24'h083)) + (({mcu[327:320], 8'b0} * 24'h0e7)) + (({mcu[335:328], 8'b0} * 24'h060)) + (({mcu[343:336], 8'b0} * -24'h060)) + (({mcu[351:344], 8'b0} * -24'h0e7)) + (({mcu[359:352], 8'b0} * -24'h0e7)) + (({mcu[367:360], 8'b0} * -24'h060)) + (({mcu[375:368], 8'b0} * 24'h060)) + (({mcu[383:376], 8'b0} * 24'h0e7)) + (({mcu[391:384], 8'b0} * 24'h02e)) + (({mcu[399:392], 8'b0} * 24'h013)) + (({mcu[407:400], 8'b0} * -24'h013)) + (({mcu[415:408], 8'b0} * -24'h02e)) + (({mcu[423:416], 8'b0} * -24'h02e)) + (({mcu[431:424], 8'b0} * -24'h013)) + (({mcu[439:432], 8'b0} * 24'h013)) + (({mcu[447:440], 8'b0} * 24'h02e)) + (({mcu[455:448], 8'b0} * -24'h0c4)) + (({mcu[463:456], 8'b0} * -24'h051)) + (({mcu[471:464], 8'b0} * 24'h051)) + (({mcu[479:472], 8'b0} * 24'h0c4)) + (({mcu[487:480], 8'b0} * 24'h0c4)) + (({mcu[495:488], 8'b0} * 24'h051)) + (({mcu[503:496], 8'b0} * -24'h051)) + (({mcu[511:504], 8'b0} * -24'h0c4));
	wire[47:0] cos33_term = (({mcu[7:0], 8'b0} * 24'h0b0)) + (({mcu[15:8], 8'b0} * -24'h029)) + (({mcu[23:16], 8'b0} * -24'h0d0)) + (({mcu[31:24], 8'b0} * -24'h076)) + (({mcu[39:32], 8'b0} * 24'h076)) + (({mcu[47:40], 8'b0} * 24'h0d0)) + (({mcu[55:48], 8'b0} * 24'h029)) + (({mcu[63:56], 8'b0} * -24'h0b0)) + (({mcu[71:64], 8'b0} * -24'h029)) + (({mcu[79:72], 8'b0} * 24'h009)) + (({mcu[87:80], 8'b0} * 24'h030)) + (({mcu[95:88], 8'b0} * 24'h01b)) + (({mcu[103:96], 8'b0} * -24'h01b)) + (({mcu[111:104], 8'b0} * -24'h030)) + (({mcu[119:112], 8'b0} * -24'h009)) + (({mcu[127:120], 8'b0} * 24'h029)) + (({mcu[135:128], 8'b0} * -24'h0d0)) + (({mcu[143:136], 8'b0} * 24'h030)) + (({mcu[151:144], 8'b0} * 24'h0f6)) + (({mcu[159:152], 8'b0} * 24'h08b)) + (({mcu[167:160], 8'b0} * -24'h08b)) + (({mcu[175:168], 8'b0} * -24'h0f6)) + (({mcu[183:176], 8'b0} * -24'h030)) + (({mcu[191:184], 8'b0} * 24'h0d0)) + (({mcu[199:192], 8'b0} * -24'h076)) + (({mcu[207:200], 8'b0} * 24'h01b)) + (({mcu[215:208], 8'b0} * 24'h08b)) + (({mcu[223:216], 8'b0} * 24'h04f)) + (({mcu[231:224], 8'b0} * -24'h04f)) + (({mcu[239:232], 8'b0} * -24'h08b)) + (({mcu[247:240], 8'b0} * -24'h01b)) + (({mcu[255:248], 8'b0} * 24'h076)) + (({mcu[263:256], 8'b0} * 24'h076)) + (({mcu[271:264], 8'b0} * -24'h01b)) + (({mcu[279:272], 8'b0} * -24'h08b)) + (({mcu[287:280], 8'b0} * -24'h04f)) + (({mcu[295:288], 8'b0} * 24'h04f)) + (({mcu[303:296], 8'b0} * 24'h08b)) + (({mcu[311:304], 8'b0} * 24'h01b)) + (({mcu[319:312], 8'b0} * -24'h076)) + (({mcu[327:320], 8'b0} * 24'h0d0)) + (({mcu[335:328], 8'b0} * -24'h030)) + (({mcu[343:336], 8'b0} * -24'h0f6)) + (({mcu[351:344], 8'b0} * -24'h08b)) + (({mcu[359:352], 8'b0} * 24'h08b)) + (({mcu[367:360], 8'b0} * 24'h0f6)) + (({mcu[375:368], 8'b0} * 24'h030)) + (({mcu[383:376], 8'b0} * -24'h0d0)) + (({mcu[391:384], 8'b0} * 24'h029)) + (({mcu[399:392], 8'b0} * -24'h009)) + (({mcu[407:400], 8'b0} * -24'h030)) + (({mcu[415:408], 8'b0} * -24'h01b)) + (({mcu[423:416], 8'b0} * 24'h01b)) + (({mcu[431:424], 8'b0} * 24'h030)) + (({mcu[439:432], 8'b0} * 24'h009)) + (({mcu[447:440], 8'b0} * -24'h029)) + (({mcu[455:448], 8'b0} * -24'h0b0)) + (({mcu[463:456], 8'b0} * 24'h029)) + (({mcu[471:464], 8'b0} * 24'h0d0)) + (({mcu[479:472], 8'b0} * 24'h076)) + (({mcu[487:480], 8'b0} * -24'h076)) + (({mcu[495:488], 8'b0} * -24'h0d0)) + (({mcu[503:496], 8'b0} * -24'h029)) + (({mcu[511:504], 8'b0} * 24'h0b0));
	wire[47:0] cos34_term = (({mcu[7:0], 8'b0} * 24'h096)) + (({mcu[15:8], 8'b0} * -24'h096)) + (({mcu[23:16], 8'b0} * -24'h096)) + (({mcu[31:24], 8'b0} * 24'h096)) + (({mcu[39:32], 8'b0} * 24'h096)) + (({mcu[47:40], 8'b0} * -24'h096)) + (({mcu[55:48], 8'b0} * -24'h096)) + (({mcu[63:56], 8'b0} * 24'h096)) + (({mcu[71:64], 8'b0} * -24'h023)) + (({mcu[79:72], 8'b0} * 24'h023)) + (({mcu[87:80], 8'b0} * 24'h023)) + (({mcu[95:88], 8'b0} * -24'h023)) + (({mcu[103:96], 8'b0} * -24'h023)) + (({mcu[111:104], 8'b0} * 24'h023)) + (({mcu[119:112], 8'b0} * 24'h023)) + (({mcu[127:120], 8'b0} * -24'h023)) + (({mcu[135:128], 8'b0} * -24'h0b1)) + (({mcu[143:136], 8'b0} * 24'h0b1)) + (({mcu[151:144], 8'b0} * 24'h0b1)) + (({mcu[159:152], 8'b0} * -24'h0b1)) + (({mcu[167:160], 8'b0} * -24'h0b1)) + (({mcu[175:168], 8'b0} * 24'h0b1)) + (({mcu[183:176], 8'b0} * 24'h0b1)) + (({mcu[191:184], 8'b0} * -24'h0b1)) + (({mcu[199:192], 8'b0} * -24'h064)) + (({mcu[207:200], 8'b0} * 24'h064)) + (({mcu[215:208], 8'b0} * 24'h064)) + (({mcu[223:216], 8'b0} * -24'h064)) + (({mcu[231:224], 8'b0} * -24'h064)) + (({mcu[239:232], 8'b0} * 24'h064)) + (({mcu[247:240], 8'b0} * 24'h064)) + (({mcu[255:248], 8'b0} * -24'h064)) + (({mcu[263:256], 8'b0} * 24'h064)) + (({mcu[271:264], 8'b0} * -24'h064)) + (({mcu[279:272], 8'b0} * -24'h064)) + (({mcu[287:280], 8'b0} * 24'h064)) + (({mcu[295:288], 8'b0} * 24'h064)) + (({mcu[303:296], 8'b0} * -24'h064)) + (({mcu[311:304], 8'b0} * -24'h064)) + (({mcu[319:312], 8'b0} * 24'h064)) + (({mcu[327:320], 8'b0} * 24'h0b1)) + (({mcu[335:328], 8'b0} * -24'h0b1)) + (({mcu[343:336], 8'b0} * -24'h0b1)) + (({mcu[351:344], 8'b0} * 24'h0b1)) + (({mcu[359:352], 8'b0} * 24'h0b1)) + (({mcu[367:360], 8'b0} * -24'h0b1)) + (({mcu[375:368], 8'b0} * -24'h0b1)) + (({mcu[383:376], 8'b0} * 24'h0b1)) + (({mcu[391:384], 8'b0} * 24'h023)) + (({mcu[399:392], 8'b0} * -24'h023)) + (({mcu[407:400], 8'b0} * -24'h023)) + (({mcu[415:408], 8'b0} * 24'h023)) + (({mcu[423:416], 8'b0} * 24'h023)) + (({mcu[431:424], 8'b0} * -24'h023)) + (({mcu[439:432], 8'b0} * -24'h023)) + (({mcu[447:440], 8'b0} * 24'h023)) + (({mcu[455:448], 8'b0} * -24'h096)) + (({mcu[463:456], 8'b0} * 24'h096)) + (({mcu[471:464], 8'b0} * 24'h096)) + (({mcu[479:472], 8'b0} * -24'h096)) + (({mcu[487:480], 8'b0} * -24'h096)) + (({mcu[495:488], 8'b0} * 24'h096)) + (({mcu[503:496], 8'b0} * 24'h096)) + (({mcu[511:504], 8'b0} * -24'h096));
	wire[47:0] cos35_term = (({mcu[7:0], 8'b0} * 24'h076)) + (({mcu[15:8], 8'b0} * -24'h0d0)) + (({mcu[23:16], 8'b0} * 24'h029)) + (({mcu[31:24], 8'b0} * 24'h0b0)) + (({mcu[39:32], 8'b0} * -24'h0b0)) + (({mcu[47:40], 8'b0} * -24'h029)) + (({mcu[55:48], 8'b0} * 24'h0d0)) + (({mcu[63:56], 8'b0} * -24'h076)) + (({mcu[71:64], 8'b0} * -24'h01b)) + (({mcu[79:72], 8'b0} * 24'h030)) + (({mcu[87:80], 8'b0} * -24'h009)) + (({mcu[95:88], 8'b0} * -24'h029)) + (({mcu[103:96], 8'b0} * 24'h029)) + (({mcu[111:104], 8'b0} * 24'h009)) + (({mcu[119:112], 8'b0} * -24'h030)) + (({mcu[127:120], 8'b0} * 24'h01b)) + (({mcu[135:128], 8'b0} * -24'h08b)) + (({mcu[143:136], 8'b0} * 24'h0f6)) + (({mcu[151:144], 8'b0} * -24'h030)) + (({mcu[159:152], 8'b0} * -24'h0d0)) + (({mcu[167:160], 8'b0} * 24'h0d0)) + (({mcu[175:168], 8'b0} * 24'h030)) + (({mcu[183:176], 8'b0} * -24'h0f6)) + (({mcu[191:184], 8'b0} * 24'h08b)) + (({mcu[199:192], 8'b0} * -24'h04f)) + (({mcu[207:200], 8'b0} * 24'h08b)) + (({mcu[215:208], 8'b0} * -24'h01b)) + (({mcu[223:216], 8'b0} * -24'h076)) + (({mcu[231:224], 8'b0} * 24'h076)) + (({mcu[239:232], 8'b0} * 24'h01b)) + (({mcu[247:240], 8'b0} * -24'h08b)) + (({mcu[255:248], 8'b0} * 24'h04f)) + (({mcu[263:256], 8'b0} * 24'h04f)) + (({mcu[271:264], 8'b0} * -24'h08b)) + (({mcu[279:272], 8'b0} * 24'h01b)) + (({mcu[287:280], 8'b0} * 24'h076)) + (({mcu[295:288], 8'b0} * -24'h076)) + (({mcu[303:296], 8'b0} * -24'h01b)) + (({mcu[311:304], 8'b0} * 24'h08b)) + (({mcu[319:312], 8'b0} * -24'h04f)) + (({mcu[327:320], 8'b0} * 24'h08b)) + (({mcu[335:328], 8'b0} * -24'h0f6)) + (({mcu[343:336], 8'b0} * 24'h030)) + (({mcu[351:344], 8'b0} * 24'h0d0)) + (({mcu[359:352], 8'b0} * -24'h0d0)) + (({mcu[367:360], 8'b0} * -24'h030)) + (({mcu[375:368], 8'b0} * 24'h0f6)) + (({mcu[383:376], 8'b0} * -24'h08b)) + (({mcu[391:384], 8'b0} * 24'h01b)) + (({mcu[399:392], 8'b0} * -24'h030)) + (({mcu[407:400], 8'b0} * 24'h009)) + (({mcu[415:408], 8'b0} * 24'h029)) + (({mcu[423:416], 8'b0} * -24'h029)) + (({mcu[431:424], 8'b0} * -24'h009)) + (({mcu[439:432], 8'b0} * 24'h030)) + (({mcu[447:440], 8'b0} * -24'h01b)) + (({mcu[455:448], 8'b0} * -24'h076)) + (({mcu[463:456], 8'b0} * 24'h0d0)) + (({mcu[471:464], 8'b0} * -24'h029)) + (({mcu[479:472], 8'b0} * -24'h0b0)) + (({mcu[487:480], 8'b0} * 24'h0b0)) + (({mcu[495:488], 8'b0} * 24'h029)) + (({mcu[503:496], 8'b0} * -24'h0d0)) + (({mcu[511:504], 8'b0} * 24'h076));
	wire[47:0] cos36_term = (({mcu[7:0], 8'b0} * 24'h051)) + (({mcu[15:8], 8'b0} * -24'h0c4)) + (({mcu[23:16], 8'b0} * 24'h0c4)) + (({mcu[31:24], 8'b0} * -24'h051)) + (({mcu[39:32], 8'b0} * -24'h051)) + (({mcu[47:40], 8'b0} * 24'h0c4)) + (({mcu[55:48], 8'b0} * -24'h0c4)) + (({mcu[63:56], 8'b0} * 24'h051)) + (({mcu[71:64], 8'b0} * -24'h013)) + (({mcu[79:72], 8'b0} * 24'h02e)) + (({mcu[87:80], 8'b0} * -24'h02e)) + (({mcu[95:88], 8'b0} * 24'h013)) + (({mcu[103:96], 8'b0} * 24'h013)) + (({mcu[111:104], 8'b0} * -24'h02e)) + (({mcu[119:112], 8'b0} * 24'h02e)) + (({mcu[127:120], 8'b0} * -24'h013)) + (({mcu[135:128], 8'b0} * -24'h060)) + (({mcu[143:136], 8'b0} * 24'h0e7)) + (({mcu[151:144], 8'b0} * -24'h0e7)) + (({mcu[159:152], 8'b0} * 24'h060)) + (({mcu[167:160], 8'b0} * 24'h060)) + (({mcu[175:168], 8'b0} * -24'h0e7)) + (({mcu[183:176], 8'b0} * 24'h0e7)) + (({mcu[191:184], 8'b0} * -24'h060)) + (({mcu[199:192], 8'b0} * -24'h036)) + (({mcu[207:200], 8'b0} * 24'h083)) + (({mcu[215:208], 8'b0} * -24'h083)) + (({mcu[223:216], 8'b0} * 24'h036)) + (({mcu[231:224], 8'b0} * 24'h036)) + (({mcu[239:232], 8'b0} * -24'h083)) + (({mcu[247:240], 8'b0} * 24'h083)) + (({mcu[255:248], 8'b0} * -24'h036)) + (({mcu[263:256], 8'b0} * 24'h036)) + (({mcu[271:264], 8'b0} * -24'h083)) + (({mcu[279:272], 8'b0} * 24'h083)) + (({mcu[287:280], 8'b0} * -24'h036)) + (({mcu[295:288], 8'b0} * -24'h036)) + (({mcu[303:296], 8'b0} * 24'h083)) + (({mcu[311:304], 8'b0} * -24'h083)) + (({mcu[319:312], 8'b0} * 24'h036)) + (({mcu[327:320], 8'b0} * 24'h060)) + (({mcu[335:328], 8'b0} * -24'h0e7)) + (({mcu[343:336], 8'b0} * 24'h0e7)) + (({mcu[351:344], 8'b0} * -24'h060)) + (({mcu[359:352], 8'b0} * -24'h060)) + (({mcu[367:360], 8'b0} * 24'h0e7)) + (({mcu[375:368], 8'b0} * -24'h0e7)) + (({mcu[383:376], 8'b0} * 24'h060)) + (({mcu[391:384], 8'b0} * 24'h013)) + (({mcu[399:392], 8'b0} * -24'h02e)) + (({mcu[407:400], 8'b0} * 24'h02e)) + (({mcu[415:408], 8'b0} * -24'h013)) + (({mcu[423:416], 8'b0} * -24'h013)) + (({mcu[431:424], 8'b0} * 24'h02e)) + (({mcu[439:432], 8'b0} * -24'h02e)) + (({mcu[447:440], 8'b0} * 24'h013)) + (({mcu[455:448], 8'b0} * -24'h051)) + (({mcu[463:456], 8'b0} * 24'h0c4)) + (({mcu[471:464], 8'b0} * -24'h0c4)) + (({mcu[479:472], 8'b0} * 24'h051)) + (({mcu[487:480], 8'b0} * 24'h051)) + (({mcu[495:488], 8'b0} * -24'h0c4)) + (({mcu[503:496], 8'b0} * 24'h0c4)) + (({mcu[511:504], 8'b0} * -24'h051));
	wire[47:0] cos37_term = (({mcu[7:0], 8'b0} * 24'h029)) + (({mcu[15:8], 8'b0} * -24'h076)) + (({mcu[23:16], 8'b0} * 24'h0b0)) + (({mcu[31:24], 8'b0} * -24'h0d0)) + (({mcu[39:32], 8'b0} * 24'h0d0)) + (({mcu[47:40], 8'b0} * -24'h0b0)) + (({mcu[55:48], 8'b0} * 24'h076)) + (({mcu[63:56], 8'b0} * -24'h029)) + (({mcu[71:64], 8'b0} * -24'h009)) + (({mcu[79:72], 8'b0} * 24'h01b)) + (({mcu[87:80], 8'b0} * -24'h029)) + (({mcu[95:88], 8'b0} * 24'h030)) + (({mcu[103:96], 8'b0} * -24'h030)) + (({mcu[111:104], 8'b0} * 24'h029)) + (({mcu[119:112], 8'b0} * -24'h01b)) + (({mcu[127:120], 8'b0} * 24'h009)) + (({mcu[135:128], 8'b0} * -24'h030)) + (({mcu[143:136], 8'b0} * 24'h08b)) + (({mcu[151:144], 8'b0} * -24'h0d0)) + (({mcu[159:152], 8'b0} * 24'h0f6)) + (({mcu[167:160], 8'b0} * -24'h0f6)) + (({mcu[175:168], 8'b0} * 24'h0d0)) + (({mcu[183:176], 8'b0} * -24'h08b)) + (({mcu[191:184], 8'b0} * 24'h030)) + (({mcu[199:192], 8'b0} * -24'h01b)) + (({mcu[207:200], 8'b0} * 24'h04f)) + (({mcu[215:208], 8'b0} * -24'h076)) + (({mcu[223:216], 8'b0} * 24'h08b)) + (({mcu[231:224], 8'b0} * -24'h08b)) + (({mcu[239:232], 8'b0} * 24'h076)) + (({mcu[247:240], 8'b0} * -24'h04f)) + (({mcu[255:248], 8'b0} * 24'h01b)) + (({mcu[263:256], 8'b0} * 24'h01b)) + (({mcu[271:264], 8'b0} * -24'h04f)) + (({mcu[279:272], 8'b0} * 24'h076)) + (({mcu[287:280], 8'b0} * -24'h08b)) + (({mcu[295:288], 8'b0} * 24'h08b)) + (({mcu[303:296], 8'b0} * -24'h076)) + (({mcu[311:304], 8'b0} * 24'h04f)) + (({mcu[319:312], 8'b0} * -24'h01b)) + (({mcu[327:320], 8'b0} * 24'h030)) + (({mcu[335:328], 8'b0} * -24'h08b)) + (({mcu[343:336], 8'b0} * 24'h0d0)) + (({mcu[351:344], 8'b0} * -24'h0f6)) + (({mcu[359:352], 8'b0} * 24'h0f6)) + (({mcu[367:360], 8'b0} * -24'h0d0)) + (({mcu[375:368], 8'b0} * 24'h08b)) + (({mcu[383:376], 8'b0} * -24'h030)) + (({mcu[391:384], 8'b0} * 24'h009)) + (({mcu[399:392], 8'b0} * -24'h01b)) + (({mcu[407:400], 8'b0} * 24'h029)) + (({mcu[415:408], 8'b0} * -24'h030)) + (({mcu[423:416], 8'b0} * 24'h030)) + (({mcu[431:424], 8'b0} * -24'h029)) + (({mcu[439:432], 8'b0} * 24'h01b)) + (({mcu[447:440], 8'b0} * -24'h009)) + (({mcu[455:448], 8'b0} * -24'h029)) + (({mcu[463:456], 8'b0} * 24'h076)) + (({mcu[471:464], 8'b0} * -24'h0b0)) + (({mcu[479:472], 8'b0} * 24'h0d0)) + (({mcu[487:480], 8'b0} * -24'h0d0)) + (({mcu[495:488], 8'b0} * 24'h0b0)) + (({mcu[503:496], 8'b0} * -24'h076)) + (({mcu[511:504], 8'b0} * 24'h029));
	wire[47:0] cos40_term = (({mcu[7:0], 8'b0} * 24'h0b4)) + (({mcu[15:8], 8'b0} * 24'h0b4)) + (({mcu[23:16], 8'b0} * 24'h0b4)) + (({mcu[31:24], 8'b0} * 24'h0b4)) + (({mcu[39:32], 8'b0} * 24'h0b4)) + (({mcu[47:40], 8'b0} * 24'h0b4)) + (({mcu[55:48], 8'b0} * 24'h0b4)) + (({mcu[63:56], 8'b0} * 24'h0b4)) + (({mcu[71:64], 8'b0} * -24'h0b4)) + (({mcu[79:72], 8'b0} * -24'h0b4)) + (({mcu[87:80], 8'b0} * -24'h0b4)) + (({mcu[95:88], 8'b0} * -24'h0b4)) + (({mcu[103:96], 8'b0} * -24'h0b4)) + (({mcu[111:104], 8'b0} * -24'h0b4)) + (({mcu[119:112], 8'b0} * -24'h0b4)) + (({mcu[127:120], 8'b0} * -24'h0b4)) + (({mcu[135:128], 8'b0} * -24'h0b4)) + (({mcu[143:136], 8'b0} * -24'h0b4)) + (({mcu[151:144], 8'b0} * -24'h0b4)) + (({mcu[159:152], 8'b0} * -24'h0b4)) + (({mcu[167:160], 8'b0} * -24'h0b4)) + (({mcu[175:168], 8'b0} * -24'h0b4)) + (({mcu[183:176], 8'b0} * -24'h0b4)) + (({mcu[191:184], 8'b0} * -24'h0b4)) + (({mcu[199:192], 8'b0} * 24'h0b4)) + (({mcu[207:200], 8'b0} * 24'h0b4)) + (({mcu[215:208], 8'b0} * 24'h0b4)) + (({mcu[223:216], 8'b0} * 24'h0b4)) + (({mcu[231:224], 8'b0} * 24'h0b4)) + (({mcu[239:232], 8'b0} * 24'h0b4)) + (({mcu[247:240], 8'b0} * 24'h0b4)) + (({mcu[255:248], 8'b0} * 24'h0b4)) + (({mcu[263:256], 8'b0} * 24'h0b4)) + (({mcu[271:264], 8'b0} * 24'h0b4)) + (({mcu[279:272], 8'b0} * 24'h0b4)) + (({mcu[287:280], 8'b0} * 24'h0b4)) + (({mcu[295:288], 8'b0} * 24'h0b4)) + (({mcu[303:296], 8'b0} * 24'h0b4)) + (({mcu[311:304], 8'b0} * 24'h0b4)) + (({mcu[319:312], 8'b0} * 24'h0b4)) + (({mcu[327:320], 8'b0} * -24'h0b4)) + (({mcu[335:328], 8'b0} * -24'h0b4)) + (({mcu[343:336], 8'b0} * -24'h0b4)) + (({mcu[351:344], 8'b0} * -24'h0b4)) + (({mcu[359:352], 8'b0} * -24'h0b4)) + (({mcu[367:360], 8'b0} * -24'h0b4)) + (({mcu[375:368], 8'b0} * -24'h0b4)) + (({mcu[383:376], 8'b0} * -24'h0b4)) + (({mcu[391:384], 8'b0} * -24'h0b4)) + (({mcu[399:392], 8'b0} * -24'h0b4)) + (({mcu[407:400], 8'b0} * -24'h0b4)) + (({mcu[415:408], 8'b0} * -24'h0b4)) + (({mcu[423:416], 8'b0} * -24'h0b4)) + (({mcu[431:424], 8'b0} * -24'h0b4)) + (({mcu[439:432], 8'b0} * -24'h0b4)) + (({mcu[447:440], 8'b0} * -24'h0b4)) + (({mcu[455:448], 8'b0} * 24'h0b4)) + (({mcu[463:456], 8'b0} * 24'h0b4)) + (({mcu[471:464], 8'b0} * 24'h0b4)) + (({mcu[479:472], 8'b0} * 24'h0b4)) + (({mcu[487:480], 8'b0} * 24'h0b4)) + (({mcu[495:488], 8'b0} * 24'h0b4)) + (({mcu[503:496], 8'b0} * 24'h0b4)) + (({mcu[511:504], 8'b0} * 24'h0b4));
	wire[47:0] cos41_term = (({mcu[7:0], 8'b0} * 24'h0b1)) + (({mcu[15:8], 8'b0} * 24'h096)) + (({mcu[23:16], 8'b0} * 24'h064)) + (({mcu[31:24], 8'b0} * 24'h023)) + (({mcu[39:32], 8'b0} * -24'h023)) + (({mcu[47:40], 8'b0} * -24'h064)) + (({mcu[55:48], 8'b0} * -24'h096)) + (({mcu[63:56], 8'b0} * -24'h0b1)) + (({mcu[71:64], 8'b0} * -24'h0b1)) + (({mcu[79:72], 8'b0} * -24'h096)) + (({mcu[87:80], 8'b0} * -24'h064)) + (({mcu[95:88], 8'b0} * -24'h023)) + (({mcu[103:96], 8'b0} * 24'h023)) + (({mcu[111:104], 8'b0} * 24'h064)) + (({mcu[119:112], 8'b0} * 24'h096)) + (({mcu[127:120], 8'b0} * 24'h0b1)) + (({mcu[135:128], 8'b0} * -24'h0b1)) + (({mcu[143:136], 8'b0} * -24'h096)) + (({mcu[151:144], 8'b0} * -24'h064)) + (({mcu[159:152], 8'b0} * -24'h023)) + (({mcu[167:160], 8'b0} * 24'h023)) + (({mcu[175:168], 8'b0} * 24'h064)) + (({mcu[183:176], 8'b0} * 24'h096)) + (({mcu[191:184], 8'b0} * 24'h0b1)) + (({mcu[199:192], 8'b0} * 24'h0b1)) + (({mcu[207:200], 8'b0} * 24'h096)) + (({mcu[215:208], 8'b0} * 24'h064)) + (({mcu[223:216], 8'b0} * 24'h023)) + (({mcu[231:224], 8'b0} * -24'h023)) + (({mcu[239:232], 8'b0} * -24'h064)) + (({mcu[247:240], 8'b0} * -24'h096)) + (({mcu[255:248], 8'b0} * -24'h0b1)) + (({mcu[263:256], 8'b0} * 24'h0b1)) + (({mcu[271:264], 8'b0} * 24'h096)) + (({mcu[279:272], 8'b0} * 24'h064)) + (({mcu[287:280], 8'b0} * 24'h023)) + (({mcu[295:288], 8'b0} * -24'h023)) + (({mcu[303:296], 8'b0} * -24'h064)) + (({mcu[311:304], 8'b0} * -24'h096)) + (({mcu[319:312], 8'b0} * -24'h0b1)) + (({mcu[327:320], 8'b0} * -24'h0b1)) + (({mcu[335:328], 8'b0} * -24'h096)) + (({mcu[343:336], 8'b0} * -24'h064)) + (({mcu[351:344], 8'b0} * -24'h023)) + (({mcu[359:352], 8'b0} * 24'h023)) + (({mcu[367:360], 8'b0} * 24'h064)) + (({mcu[375:368], 8'b0} * 24'h096)) + (({mcu[383:376], 8'b0} * 24'h0b1)) + (({mcu[391:384], 8'b0} * -24'h0b1)) + (({mcu[399:392], 8'b0} * -24'h096)) + (({mcu[407:400], 8'b0} * -24'h064)) + (({mcu[415:408], 8'b0} * -24'h023)) + (({mcu[423:416], 8'b0} * 24'h023)) + (({mcu[431:424], 8'b0} * 24'h064)) + (({mcu[439:432], 8'b0} * 24'h096)) + (({mcu[447:440], 8'b0} * 24'h0b1)) + (({mcu[455:448], 8'b0} * 24'h0b1)) + (({mcu[463:456], 8'b0} * 24'h096)) + (({mcu[471:464], 8'b0} * 24'h064)) + (({mcu[479:472], 8'b0} * 24'h023)) + (({mcu[487:480], 8'b0} * -24'h023)) + (({mcu[495:488], 8'b0} * -24'h064)) + (({mcu[503:496], 8'b0} * -24'h096)) + (({mcu[511:504], 8'b0} * -24'h0b1));
	wire[47:0] cos42_term = (({mcu[7:0], 8'b0} * 24'h0a7)) + (({mcu[15:8], 8'b0} * 24'h045)) + (({mcu[23:16], 8'b0} * -24'h045)) + (({mcu[31:24], 8'b0} * -24'h0a7)) + (({mcu[39:32], 8'b0} * -24'h0a7)) + (({mcu[47:40], 8'b0} * -24'h045)) + (({mcu[55:48], 8'b0} * 24'h045)) + (({mcu[63:56], 8'b0} * 24'h0a7)) + (({mcu[71:64], 8'b0} * -24'h0a7)) + (({mcu[79:72], 8'b0} * -24'h045)) + (({mcu[87:80], 8'b0} * 24'h045)) + (({mcu[95:88], 8'b0} * 24'h0a7)) + (({mcu[103:96], 8'b0} * 24'h0a7)) + (({mcu[111:104], 8'b0} * 24'h045)) + (({mcu[119:112], 8'b0} * -24'h045)) + (({mcu[127:120], 8'b0} * -24'h0a7)) + (({mcu[135:128], 8'b0} * -24'h0a7)) + (({mcu[143:136], 8'b0} * -24'h045)) + (({mcu[151:144], 8'b0} * 24'h045)) + (({mcu[159:152], 8'b0} * 24'h0a7)) + (({mcu[167:160], 8'b0} * 24'h0a7)) + (({mcu[175:168], 8'b0} * 24'h045)) + (({mcu[183:176], 8'b0} * -24'h045)) + (({mcu[191:184], 8'b0} * -24'h0a7)) + (({mcu[199:192], 8'b0} * 24'h0a7)) + (({mcu[207:200], 8'b0} * 24'h045)) + (({mcu[215:208], 8'b0} * -24'h045)) + (({mcu[223:216], 8'b0} * -24'h0a7)) + (({mcu[231:224], 8'b0} * -24'h0a7)) + (({mcu[239:232], 8'b0} * -24'h045)) + (({mcu[247:240], 8'b0} * 24'h045)) + (({mcu[255:248], 8'b0} * 24'h0a7)) + (({mcu[263:256], 8'b0} * 24'h0a7)) + (({mcu[271:264], 8'b0} * 24'h045)) + (({mcu[279:272], 8'b0} * -24'h045)) + (({mcu[287:280], 8'b0} * -24'h0a7)) + (({mcu[295:288], 8'b0} * -24'h0a7)) + (({mcu[303:296], 8'b0} * -24'h045)) + (({mcu[311:304], 8'b0} * 24'h045)) + (({mcu[319:312], 8'b0} * 24'h0a7)) + (({mcu[327:320], 8'b0} * -24'h0a7)) + (({mcu[335:328], 8'b0} * -24'h045)) + (({mcu[343:336], 8'b0} * 24'h045)) + (({mcu[351:344], 8'b0} * 24'h0a7)) + (({mcu[359:352], 8'b0} * 24'h0a7)) + (({mcu[367:360], 8'b0} * 24'h045)) + (({mcu[375:368], 8'b0} * -24'h045)) + (({mcu[383:376], 8'b0} * -24'h0a7)) + (({mcu[391:384], 8'b0} * -24'h0a7)) + (({mcu[399:392], 8'b0} * -24'h045)) + (({mcu[407:400], 8'b0} * 24'h045)) + (({mcu[415:408], 8'b0} * 24'h0a7)) + (({mcu[423:416], 8'b0} * 24'h0a7)) + (({mcu[431:424], 8'b0} * 24'h045)) + (({mcu[439:432], 8'b0} * -24'h045)) + (({mcu[447:440], 8'b0} * -24'h0a7)) + (({mcu[455:448], 8'b0} * 24'h0a7)) + (({mcu[463:456], 8'b0} * 24'h045)) + (({mcu[471:464], 8'b0} * -24'h045)) + (({mcu[479:472], 8'b0} * -24'h0a7)) + (({mcu[487:480], 8'b0} * -24'h0a7)) + (({mcu[495:488], 8'b0} * -24'h045)) + (({mcu[503:496], 8'b0} * 24'h045)) + (({mcu[511:504], 8'b0} * 24'h0a7));
	wire[47:0] cos43_term = (({mcu[7:0], 8'b0} * 24'h096)) + (({mcu[15:8], 8'b0} * -24'h023)) + (({mcu[23:16], 8'b0} * -24'h0b1)) + (({mcu[31:24], 8'b0} * -24'h064)) + (({mcu[39:32], 8'b0} * 24'h064)) + (({mcu[47:40], 8'b0} * 24'h0b1)) + (({mcu[55:48], 8'b0} * 24'h023)) + (({mcu[63:56], 8'b0} * -24'h096)) + (({mcu[71:64], 8'b0} * -24'h096)) + (({mcu[79:72], 8'b0} * 24'h023)) + (({mcu[87:80], 8'b0} * 24'h0b1)) + (({mcu[95:88], 8'b0} * 24'h064)) + (({mcu[103:96], 8'b0} * -24'h064)) + (({mcu[111:104], 8'b0} * -24'h0b1)) + (({mcu[119:112], 8'b0} * -24'h023)) + (({mcu[127:120], 8'b0} * 24'h096)) + (({mcu[135:128], 8'b0} * -24'h096)) + (({mcu[143:136], 8'b0} * 24'h023)) + (({mcu[151:144], 8'b0} * 24'h0b1)) + (({mcu[159:152], 8'b0} * 24'h064)) + (({mcu[167:160], 8'b0} * -24'h064)) + (({mcu[175:168], 8'b0} * -24'h0b1)) + (({mcu[183:176], 8'b0} * -24'h023)) + (({mcu[191:184], 8'b0} * 24'h096)) + (({mcu[199:192], 8'b0} * 24'h096)) + (({mcu[207:200], 8'b0} * -24'h023)) + (({mcu[215:208], 8'b0} * -24'h0b1)) + (({mcu[223:216], 8'b0} * -24'h064)) + (({mcu[231:224], 8'b0} * 24'h064)) + (({mcu[239:232], 8'b0} * 24'h0b1)) + (({mcu[247:240], 8'b0} * 24'h023)) + (({mcu[255:248], 8'b0} * -24'h096)) + (({mcu[263:256], 8'b0} * 24'h096)) + (({mcu[271:264], 8'b0} * -24'h023)) + (({mcu[279:272], 8'b0} * -24'h0b1)) + (({mcu[287:280], 8'b0} * -24'h064)) + (({mcu[295:288], 8'b0} * 24'h064)) + (({mcu[303:296], 8'b0} * 24'h0b1)) + (({mcu[311:304], 8'b0} * 24'h023)) + (({mcu[319:312], 8'b0} * -24'h096)) + (({mcu[327:320], 8'b0} * -24'h096)) + (({mcu[335:328], 8'b0} * 24'h023)) + (({mcu[343:336], 8'b0} * 24'h0b1)) + (({mcu[351:344], 8'b0} * 24'h064)) + (({mcu[359:352], 8'b0} * -24'h064)) + (({mcu[367:360], 8'b0} * -24'h0b1)) + (({mcu[375:368], 8'b0} * -24'h023)) + (({mcu[383:376], 8'b0} * 24'h096)) + (({mcu[391:384], 8'b0} * -24'h096)) + (({mcu[399:392], 8'b0} * 24'h023)) + (({mcu[407:400], 8'b0} * 24'h0b1)) + (({mcu[415:408], 8'b0} * 24'h064)) + (({mcu[423:416], 8'b0} * -24'h064)) + (({mcu[431:424], 8'b0} * -24'h0b1)) + (({mcu[439:432], 8'b0} * -24'h023)) + (({mcu[447:440], 8'b0} * 24'h096)) + (({mcu[455:448], 8'b0} * 24'h096)) + (({mcu[463:456], 8'b0} * -24'h023)) + (({mcu[471:464], 8'b0} * -24'h0b1)) + (({mcu[479:472], 8'b0} * -24'h064)) + (({mcu[487:480], 8'b0} * 24'h064)) + (({mcu[495:488], 8'b0} * 24'h0b1)) + (({mcu[503:496], 8'b0} * 24'h023)) + (({mcu[511:504], 8'b0} * -24'h096));
	wire[47:0] cos44_term = (({mcu[7:0], 8'b0} * 24'h080)) + (({mcu[15:8], 8'b0} * -24'h080)) + (({mcu[23:16], 8'b0} * -24'h080)) + (({mcu[31:24], 8'b0} * 24'h080)) + (({mcu[39:32], 8'b0} * 24'h080)) + (({mcu[47:40], 8'b0} * -24'h080)) + (({mcu[55:48], 8'b0} * -24'h080)) + (({mcu[63:56], 8'b0} * 24'h080)) + (({mcu[71:64], 8'b0} * -24'h080)) + (({mcu[79:72], 8'b0} * 24'h080)) + (({mcu[87:80], 8'b0} * 24'h080)) + (({mcu[95:88], 8'b0} * -24'h080)) + (({mcu[103:96], 8'b0} * -24'h080)) + (({mcu[111:104], 8'b0} * 24'h080)) + (({mcu[119:112], 8'b0} * 24'h080)) + (({mcu[127:120], 8'b0} * -24'h080)) + (({mcu[135:128], 8'b0} * -24'h080)) + (({mcu[143:136], 8'b0} * 24'h080)) + (({mcu[151:144], 8'b0} * 24'h080)) + (({mcu[159:152], 8'b0} * -24'h080)) + (({mcu[167:160], 8'b0} * -24'h080)) + (({mcu[175:168], 8'b0} * 24'h080)) + (({mcu[183:176], 8'b0} * 24'h080)) + (({mcu[191:184], 8'b0} * -24'h080)) + (({mcu[199:192], 8'b0} * 24'h080)) + (({mcu[207:200], 8'b0} * -24'h080)) + (({mcu[215:208], 8'b0} * -24'h080)) + (({mcu[223:216], 8'b0} * 24'h080)) + (({mcu[231:224], 8'b0} * 24'h080)) + (({mcu[239:232], 8'b0} * -24'h080)) + (({mcu[247:240], 8'b0} * -24'h080)) + (({mcu[255:248], 8'b0} * 24'h080)) + (({mcu[263:256], 8'b0} * 24'h080)) + (({mcu[271:264], 8'b0} * -24'h080)) + (({mcu[279:272], 8'b0} * -24'h080)) + (({mcu[287:280], 8'b0} * 24'h080)) + (({mcu[295:288], 8'b0} * 24'h080)) + (({mcu[303:296], 8'b0} * -24'h080)) + (({mcu[311:304], 8'b0} * -24'h080)) + (({mcu[319:312], 8'b0} * 24'h080)) + (({mcu[327:320], 8'b0} * -24'h080)) + (({mcu[335:328], 8'b0} * 24'h080)) + (({mcu[343:336], 8'b0} * 24'h080)) + (({mcu[351:344], 8'b0} * -24'h080)) + (({mcu[359:352], 8'b0} * -24'h080)) + (({mcu[367:360], 8'b0} * 24'h080)) + (({mcu[375:368], 8'b0} * 24'h080)) + (({mcu[383:376], 8'b0} * -24'h080)) + (({mcu[391:384], 8'b0} * -24'h080)) + (({mcu[399:392], 8'b0} * 24'h080)) + (({mcu[407:400], 8'b0} * 24'h080)) + (({mcu[415:408], 8'b0} * -24'h080)) + (({mcu[423:416], 8'b0} * -24'h080)) + (({mcu[431:424], 8'b0} * 24'h080)) + (({mcu[439:432], 8'b0} * 24'h080)) + (({mcu[447:440], 8'b0} * -24'h080)) + (({mcu[455:448], 8'b0} * 24'h080)) + (({mcu[463:456], 8'b0} * -24'h080)) + (({mcu[471:464], 8'b0} * -24'h080)) + (({mcu[479:472], 8'b0} * 24'h080)) + (({mcu[487:480], 8'b0} * 24'h080)) + (({mcu[495:488], 8'b0} * -24'h080)) + (({mcu[503:496], 8'b0} * -24'h080)) + (({mcu[511:504], 8'b0} * 24'h080));
	wire[47:0] cos45_term = (({mcu[7:0], 8'b0} * 24'h064)) + (({mcu[15:8], 8'b0} * -24'h0b1)) + (({mcu[23:16], 8'b0} * 24'h023)) + (({mcu[31:24], 8'b0} * 24'h096)) + (({mcu[39:32], 8'b0} * -24'h096)) + (({mcu[47:40], 8'b0} * -24'h023)) + (({mcu[55:48], 8'b0} * 24'h0b1)) + (({mcu[63:56], 8'b0} * -24'h064)) + (({mcu[71:64], 8'b0} * -24'h064)) + (({mcu[79:72], 8'b0} * 24'h0b1)) + (({mcu[87:80], 8'b0} * -24'h023)) + (({mcu[95:88], 8'b0} * -24'h096)) + (({mcu[103:96], 8'b0} * 24'h096)) + (({mcu[111:104], 8'b0} * 24'h023)) + (({mcu[119:112], 8'b0} * -24'h0b1)) + (({mcu[127:120], 8'b0} * 24'h064)) + (({mcu[135:128], 8'b0} * -24'h064)) + (({mcu[143:136], 8'b0} * 24'h0b1)) + (({mcu[151:144], 8'b0} * -24'h023)) + (({mcu[159:152], 8'b0} * -24'h096)) + (({mcu[167:160], 8'b0} * 24'h096)) + (({mcu[175:168], 8'b0} * 24'h023)) + (({mcu[183:176], 8'b0} * -24'h0b1)) + (({mcu[191:184], 8'b0} * 24'h064)) + (({mcu[199:192], 8'b0} * 24'h064)) + (({mcu[207:200], 8'b0} * -24'h0b1)) + (({mcu[215:208], 8'b0} * 24'h023)) + (({mcu[223:216], 8'b0} * 24'h096)) + (({mcu[231:224], 8'b0} * -24'h096)) + (({mcu[239:232], 8'b0} * -24'h023)) + (({mcu[247:240], 8'b0} * 24'h0b1)) + (({mcu[255:248], 8'b0} * -24'h064)) + (({mcu[263:256], 8'b0} * 24'h064)) + (({mcu[271:264], 8'b0} * -24'h0b1)) + (({mcu[279:272], 8'b0} * 24'h023)) + (({mcu[287:280], 8'b0} * 24'h096)) + (({mcu[295:288], 8'b0} * -24'h096)) + (({mcu[303:296], 8'b0} * -24'h023)) + (({mcu[311:304], 8'b0} * 24'h0b1)) + (({mcu[319:312], 8'b0} * -24'h064)) + (({mcu[327:320], 8'b0} * -24'h064)) + (({mcu[335:328], 8'b0} * 24'h0b1)) + (({mcu[343:336], 8'b0} * -24'h023)) + (({mcu[351:344], 8'b0} * -24'h096)) + (({mcu[359:352], 8'b0} * 24'h096)) + (({mcu[367:360], 8'b0} * 24'h023)) + (({mcu[375:368], 8'b0} * -24'h0b1)) + (({mcu[383:376], 8'b0} * 24'h064)) + (({mcu[391:384], 8'b0} * -24'h064)) + (({mcu[399:392], 8'b0} * 24'h0b1)) + (({mcu[407:400], 8'b0} * -24'h023)) + (({mcu[415:408], 8'b0} * -24'h096)) + (({mcu[423:416], 8'b0} * 24'h096)) + (({mcu[431:424], 8'b0} * 24'h023)) + (({mcu[439:432], 8'b0} * -24'h0b1)) + (({mcu[447:440], 8'b0} * 24'h064)) + (({mcu[455:448], 8'b0} * 24'h064)) + (({mcu[463:456], 8'b0} * -24'h0b1)) + (({mcu[471:464], 8'b0} * 24'h023)) + (({mcu[479:472], 8'b0} * 24'h096)) + (({mcu[487:480], 8'b0} * -24'h096)) + (({mcu[495:488], 8'b0} * -24'h023)) + (({mcu[503:496], 8'b0} * 24'h0b1)) + (({mcu[511:504], 8'b0} * -24'h064));
	wire[47:0] cos46_term = (({mcu[7:0], 8'b0} * 24'h045)) + (({mcu[15:8], 8'b0} * -24'h0a7)) + (({mcu[23:16], 8'b0} * 24'h0a7)) + (({mcu[31:24], 8'b0} * -24'h045)) + (({mcu[39:32], 8'b0} * -24'h045)) + (({mcu[47:40], 8'b0} * 24'h0a7)) + (({mcu[55:48], 8'b0} * -24'h0a7)) + (({mcu[63:56], 8'b0} * 24'h045)) + (({mcu[71:64], 8'b0} * -24'h045)) + (({mcu[79:72], 8'b0} * 24'h0a7)) + (({mcu[87:80], 8'b0} * -24'h0a7)) + (({mcu[95:88], 8'b0} * 24'h045)) + (({mcu[103:96], 8'b0} * 24'h045)) + (({mcu[111:104], 8'b0} * -24'h0a7)) + (({mcu[119:112], 8'b0} * 24'h0a7)) + (({mcu[127:120], 8'b0} * -24'h045)) + (({mcu[135:128], 8'b0} * -24'h045)) + (({mcu[143:136], 8'b0} * 24'h0a7)) + (({mcu[151:144], 8'b0} * -24'h0a7)) + (({mcu[159:152], 8'b0} * 24'h045)) + (({mcu[167:160], 8'b0} * 24'h045)) + (({mcu[175:168], 8'b0} * -24'h0a7)) + (({mcu[183:176], 8'b0} * 24'h0a7)) + (({mcu[191:184], 8'b0} * -24'h045)) + (({mcu[199:192], 8'b0} * 24'h045)) + (({mcu[207:200], 8'b0} * -24'h0a7)) + (({mcu[215:208], 8'b0} * 24'h0a7)) + (({mcu[223:216], 8'b0} * -24'h045)) + (({mcu[231:224], 8'b0} * -24'h045)) + (({mcu[239:232], 8'b0} * 24'h0a7)) + (({mcu[247:240], 8'b0} * -24'h0a7)) + (({mcu[255:248], 8'b0} * 24'h045)) + (({mcu[263:256], 8'b0} * 24'h045)) + (({mcu[271:264], 8'b0} * -24'h0a7)) + (({mcu[279:272], 8'b0} * 24'h0a7)) + (({mcu[287:280], 8'b0} * -24'h045)) + (({mcu[295:288], 8'b0} * -24'h045)) + (({mcu[303:296], 8'b0} * 24'h0a7)) + (({mcu[311:304], 8'b0} * -24'h0a7)) + (({mcu[319:312], 8'b0} * 24'h045)) + (({mcu[327:320], 8'b0} * -24'h045)) + (({mcu[335:328], 8'b0} * 24'h0a7)) + (({mcu[343:336], 8'b0} * -24'h0a7)) + (({mcu[351:344], 8'b0} * 24'h045)) + (({mcu[359:352], 8'b0} * 24'h045)) + (({mcu[367:360], 8'b0} * -24'h0a7)) + (({mcu[375:368], 8'b0} * 24'h0a7)) + (({mcu[383:376], 8'b0} * -24'h045)) + (({mcu[391:384], 8'b0} * -24'h045)) + (({mcu[399:392], 8'b0} * 24'h0a7)) + (({mcu[407:400], 8'b0} * -24'h0a7)) + (({mcu[415:408], 8'b0} * 24'h045)) + (({mcu[423:416], 8'b0} * 24'h045)) + (({mcu[431:424], 8'b0} * -24'h0a7)) + (({mcu[439:432], 8'b0} * 24'h0a7)) + (({mcu[447:440], 8'b0} * -24'h045)) + (({mcu[455:448], 8'b0} * 24'h045)) + (({mcu[463:456], 8'b0} * -24'h0a7)) + (({mcu[471:464], 8'b0} * 24'h0a7)) + (({mcu[479:472], 8'b0} * -24'h045)) + (({mcu[487:480], 8'b0} * -24'h045)) + (({mcu[495:488], 8'b0} * 24'h0a7)) + (({mcu[503:496], 8'b0} * -24'h0a7)) + (({mcu[511:504], 8'b0} * 24'h045));
	wire[47:0] cos47_term = (({mcu[7:0], 8'b0} * 24'h023)) + (({mcu[15:8], 8'b0} * -24'h064)) + (({mcu[23:16], 8'b0} * 24'h096)) + (({mcu[31:24], 8'b0} * -24'h0b1)) + (({mcu[39:32], 8'b0} * 24'h0b1)) + (({mcu[47:40], 8'b0} * -24'h096)) + (({mcu[55:48], 8'b0} * 24'h064)) + (({mcu[63:56], 8'b0} * -24'h023)) + (({mcu[71:64], 8'b0} * -24'h023)) + (({mcu[79:72], 8'b0} * 24'h064)) + (({mcu[87:80], 8'b0} * -24'h096)) + (({mcu[95:88], 8'b0} * 24'h0b1)) + (({mcu[103:96], 8'b0} * -24'h0b1)) + (({mcu[111:104], 8'b0} * 24'h096)) + (({mcu[119:112], 8'b0} * -24'h064)) + (({mcu[127:120], 8'b0} * 24'h023)) + (({mcu[135:128], 8'b0} * -24'h023)) + (({mcu[143:136], 8'b0} * 24'h064)) + (({mcu[151:144], 8'b0} * -24'h096)) + (({mcu[159:152], 8'b0} * 24'h0b1)) + (({mcu[167:160], 8'b0} * -24'h0b1)) + (({mcu[175:168], 8'b0} * 24'h096)) + (({mcu[183:176], 8'b0} * -24'h064)) + (({mcu[191:184], 8'b0} * 24'h023)) + (({mcu[199:192], 8'b0} * 24'h023)) + (({mcu[207:200], 8'b0} * -24'h064)) + (({mcu[215:208], 8'b0} * 24'h096)) + (({mcu[223:216], 8'b0} * -24'h0b1)) + (({mcu[231:224], 8'b0} * 24'h0b1)) + (({mcu[239:232], 8'b0} * -24'h096)) + (({mcu[247:240], 8'b0} * 24'h064)) + (({mcu[255:248], 8'b0} * -24'h023)) + (({mcu[263:256], 8'b0} * 24'h023)) + (({mcu[271:264], 8'b0} * -24'h064)) + (({mcu[279:272], 8'b0} * 24'h096)) + (({mcu[287:280], 8'b0} * -24'h0b1)) + (({mcu[295:288], 8'b0} * 24'h0b1)) + (({mcu[303:296], 8'b0} * -24'h096)) + (({mcu[311:304], 8'b0} * 24'h064)) + (({mcu[319:312], 8'b0} * -24'h023)) + (({mcu[327:320], 8'b0} * -24'h023)) + (({mcu[335:328], 8'b0} * 24'h064)) + (({mcu[343:336], 8'b0} * -24'h096)) + (({mcu[351:344], 8'b0} * 24'h0b1)) + (({mcu[359:352], 8'b0} * -24'h0b1)) + (({mcu[367:360], 8'b0} * 24'h096)) + (({mcu[375:368], 8'b0} * -24'h064)) + (({mcu[383:376], 8'b0} * 24'h023)) + (({mcu[391:384], 8'b0} * -24'h023)) + (({mcu[399:392], 8'b0} * 24'h064)) + (({mcu[407:400], 8'b0} * -24'h096)) + (({mcu[415:408], 8'b0} * 24'h0b1)) + (({mcu[423:416], 8'b0} * -24'h0b1)) + (({mcu[431:424], 8'b0} * 24'h096)) + (({mcu[439:432], 8'b0} * -24'h064)) + (({mcu[447:440], 8'b0} * 24'h023)) + (({mcu[455:448], 8'b0} * 24'h023)) + (({mcu[463:456], 8'b0} * -24'h064)) + (({mcu[471:464], 8'b0} * 24'h096)) + (({mcu[479:472], 8'b0} * -24'h0b1)) + (({mcu[487:480], 8'b0} * 24'h0b1)) + (({mcu[495:488], 8'b0} * -24'h096)) + (({mcu[503:496], 8'b0} * 24'h064)) + (({mcu[511:504], 8'b0} * -24'h023));
	wire[47:0] cos50_term = (({mcu[7:0], 8'b0} * 24'h08e)) + (({mcu[15:8], 8'b0} * 24'h08e)) + (({mcu[23:16], 8'b0} * 24'h08e)) + (({mcu[31:24], 8'b0} * 24'h08e)) + (({mcu[39:32], 8'b0} * 24'h08e)) + (({mcu[47:40], 8'b0} * 24'h08e)) + (({mcu[55:48], 8'b0} * 24'h08e)) + (({mcu[63:56], 8'b0} * 24'h08e)) + (({mcu[71:64], 8'b0} * -24'h0fb)) + (({mcu[79:72], 8'b0} * -24'h0fb)) + (({mcu[87:80], 8'b0} * -24'h0fb)) + (({mcu[95:88], 8'b0} * -24'h0fb)) + (({mcu[103:96], 8'b0} * -24'h0fb)) + (({mcu[111:104], 8'b0} * -24'h0fb)) + (({mcu[119:112], 8'b0} * -24'h0fb)) + (({mcu[127:120], 8'b0} * -24'h0fb)) + (({mcu[135:128], 8'b0} * 24'h031)) + (({mcu[143:136], 8'b0} * 24'h031)) + (({mcu[151:144], 8'b0} * 24'h031)) + (({mcu[159:152], 8'b0} * 24'h031)) + (({mcu[167:160], 8'b0} * 24'h031)) + (({mcu[175:168], 8'b0} * 24'h031)) + (({mcu[183:176], 8'b0} * 24'h031)) + (({mcu[191:184], 8'b0} * 24'h031)) + (({mcu[199:192], 8'b0} * 24'h0d4)) + (({mcu[207:200], 8'b0} * 24'h0d4)) + (({mcu[215:208], 8'b0} * 24'h0d4)) + (({mcu[223:216], 8'b0} * 24'h0d4)) + (({mcu[231:224], 8'b0} * 24'h0d4)) + (({mcu[239:232], 8'b0} * 24'h0d4)) + (({mcu[247:240], 8'b0} * 24'h0d4)) + (({mcu[255:248], 8'b0} * 24'h0d4)) + (({mcu[263:256], 8'b0} * -24'h0d4)) + (({mcu[271:264], 8'b0} * -24'h0d4)) + (({mcu[279:272], 8'b0} * -24'h0d4)) + (({mcu[287:280], 8'b0} * -24'h0d4)) + (({mcu[295:288], 8'b0} * -24'h0d4)) + (({mcu[303:296], 8'b0} * -24'h0d4)) + (({mcu[311:304], 8'b0} * -24'h0d4)) + (({mcu[319:312], 8'b0} * -24'h0d4)) + (({mcu[327:320], 8'b0} * -24'h031)) + (({mcu[335:328], 8'b0} * -24'h031)) + (({mcu[343:336], 8'b0} * -24'h031)) + (({mcu[351:344], 8'b0} * -24'h031)) + (({mcu[359:352], 8'b0} * -24'h031)) + (({mcu[367:360], 8'b0} * -24'h031)) + (({mcu[375:368], 8'b0} * -24'h031)) + (({mcu[383:376], 8'b0} * -24'h031)) + (({mcu[391:384], 8'b0} * 24'h0fb)) + (({mcu[399:392], 8'b0} * 24'h0fb)) + (({mcu[407:400], 8'b0} * 24'h0fb)) + (({mcu[415:408], 8'b0} * 24'h0fb)) + (({mcu[423:416], 8'b0} * 24'h0fb)) + (({mcu[431:424], 8'b0} * 24'h0fb)) + (({mcu[439:432], 8'b0} * 24'h0fb)) + (({mcu[447:440], 8'b0} * 24'h0fb)) + (({mcu[455:448], 8'b0} * -24'h08e)) + (({mcu[463:456], 8'b0} * -24'h08e)) + (({mcu[471:464], 8'b0} * -24'h08e)) + (({mcu[479:472], 8'b0} * -24'h08e)) + (({mcu[487:480], 8'b0} * -24'h08e)) + (({mcu[495:488], 8'b0} * -24'h08e)) + (({mcu[503:496], 8'b0} * -24'h08e)) + (({mcu[511:504], 8'b0} * -24'h08e));
	wire[47:0] cos51_term = (({mcu[7:0], 8'b0} * 24'h08b)) + (({mcu[15:8], 8'b0} * 24'h076)) + (({mcu[23:16], 8'b0} * 24'h04f)) + (({mcu[31:24], 8'b0} * 24'h01b)) + (({mcu[39:32], 8'b0} * -24'h01b)) + (({mcu[47:40], 8'b0} * -24'h04f)) + (({mcu[55:48], 8'b0} * -24'h076)) + (({mcu[63:56], 8'b0} * -24'h08b)) + (({mcu[71:64], 8'b0} * -24'h0f6)) + (({mcu[79:72], 8'b0} * -24'h0d0)) + (({mcu[87:80], 8'b0} * -24'h08b)) + (({mcu[95:88], 8'b0} * -24'h030)) + (({mcu[103:96], 8'b0} * 24'h030)) + (({mcu[111:104], 8'b0} * 24'h08b)) + (({mcu[119:112], 8'b0} * 24'h0d0)) + (({mcu[127:120], 8'b0} * 24'h0f6)) + (({mcu[135:128], 8'b0} * 24'h030)) + (({mcu[143:136], 8'b0} * 24'h029)) + (({mcu[151:144], 8'b0} * 24'h01b)) + (({mcu[159:152], 8'b0} * 24'h009)) + (({mcu[167:160], 8'b0} * -24'h009)) + (({mcu[175:168], 8'b0} * -24'h01b)) + (({mcu[183:176], 8'b0} * -24'h029)) + (({mcu[191:184], 8'b0} * -24'h030)) + (({mcu[199:192], 8'b0} * 24'h0d0)) + (({mcu[207:200], 8'b0} * 24'h0b0)) + (({mcu[215:208], 8'b0} * 24'h076)) + (({mcu[223:216], 8'b0} * 24'h029)) + (({mcu[231:224], 8'b0} * -24'h029)) + (({mcu[239:232], 8'b0} * -24'h076)) + (({mcu[247:240], 8'b0} * -24'h0b0)) + (({mcu[255:248], 8'b0} * -24'h0d0)) + (({mcu[263:256], 8'b0} * -24'h0d0)) + (({mcu[271:264], 8'b0} * -24'h0b0)) + (({mcu[279:272], 8'b0} * -24'h076)) + (({mcu[287:280], 8'b0} * -24'h029)) + (({mcu[295:288], 8'b0} * 24'h029)) + (({mcu[303:296], 8'b0} * 24'h076)) + (({mcu[311:304], 8'b0} * 24'h0b0)) + (({mcu[319:312], 8'b0} * 24'h0d0)) + (({mcu[327:320], 8'b0} * -24'h030)) + (({mcu[335:328], 8'b0} * -24'h029)) + (({mcu[343:336], 8'b0} * -24'h01b)) + (({mcu[351:344], 8'b0} * -24'h009)) + (({mcu[359:352], 8'b0} * 24'h009)) + (({mcu[367:360], 8'b0} * 24'h01b)) + (({mcu[375:368], 8'b0} * 24'h029)) + (({mcu[383:376], 8'b0} * 24'h030)) + (({mcu[391:384], 8'b0} * 24'h0f6)) + (({mcu[399:392], 8'b0} * 24'h0d0)) + (({mcu[407:400], 8'b0} * 24'h08b)) + (({mcu[415:408], 8'b0} * 24'h030)) + (({mcu[423:416], 8'b0} * -24'h030)) + (({mcu[431:424], 8'b0} * -24'h08b)) + (({mcu[439:432], 8'b0} * -24'h0d0)) + (({mcu[447:440], 8'b0} * -24'h0f6)) + (({mcu[455:448], 8'b0} * -24'h08b)) + (({mcu[463:456], 8'b0} * -24'h076)) + (({mcu[471:464], 8'b0} * -24'h04f)) + (({mcu[479:472], 8'b0} * -24'h01b)) + (({mcu[487:480], 8'b0} * 24'h01b)) + (({mcu[495:488], 8'b0} * 24'h04f)) + (({mcu[503:496], 8'b0} * 24'h076)) + (({mcu[511:504], 8'b0} * 24'h08b));
	wire[47:0] cos52_term = (({mcu[7:0], 8'b0} * 24'h083)) + (({mcu[15:8], 8'b0} * 24'h036)) + (({mcu[23:16], 8'b0} * -24'h036)) + (({mcu[31:24], 8'b0} * -24'h083)) + (({mcu[39:32], 8'b0} * -24'h083)) + (({mcu[47:40], 8'b0} * -24'h036)) + (({mcu[55:48], 8'b0} * 24'h036)) + (({mcu[63:56], 8'b0} * 24'h083)) + (({mcu[71:64], 8'b0} * -24'h0e7)) + (({mcu[79:72], 8'b0} * -24'h060)) + (({mcu[87:80], 8'b0} * 24'h060)) + (({mcu[95:88], 8'b0} * 24'h0e7)) + (({mcu[103:96], 8'b0} * 24'h0e7)) + (({mcu[111:104], 8'b0} * 24'h060)) + (({mcu[119:112], 8'b0} * -24'h060)) + (({mcu[127:120], 8'b0} * -24'h0e7)) + (({mcu[135:128], 8'b0} * 24'h02e)) + (({mcu[143:136], 8'b0} * 24'h013)) + (({mcu[151:144], 8'b0} * -24'h013)) + (({mcu[159:152], 8'b0} * -24'h02e)) + (({mcu[167:160], 8'b0} * -24'h02e)) + (({mcu[175:168], 8'b0} * -24'h013)) + (({mcu[183:176], 8'b0} * 24'h013)) + (({mcu[191:184], 8'b0} * 24'h02e)) + (({mcu[199:192], 8'b0} * 24'h0c4)) + (({mcu[207:200], 8'b0} * 24'h051)) + (({mcu[215:208], 8'b0} * -24'h051)) + (({mcu[223:216], 8'b0} * -24'h0c4)) + (({mcu[231:224], 8'b0} * -24'h0c4)) + (({mcu[239:232], 8'b0} * -24'h051)) + (({mcu[247:240], 8'b0} * 24'h051)) + (({mcu[255:248], 8'b0} * 24'h0c4)) + (({mcu[263:256], 8'b0} * -24'h0c4)) + (({mcu[271:264], 8'b0} * -24'h051)) + (({mcu[279:272], 8'b0} * 24'h051)) + (({mcu[287:280], 8'b0} * 24'h0c4)) + (({mcu[295:288], 8'b0} * 24'h0c4)) + (({mcu[303:296], 8'b0} * 24'h051)) + (({mcu[311:304], 8'b0} * -24'h051)) + (({mcu[319:312], 8'b0} * -24'h0c4)) + (({mcu[327:320], 8'b0} * -24'h02e)) + (({mcu[335:328], 8'b0} * -24'h013)) + (({mcu[343:336], 8'b0} * 24'h013)) + (({mcu[351:344], 8'b0} * 24'h02e)) + (({mcu[359:352], 8'b0} * 24'h02e)) + (({mcu[367:360], 8'b0} * 24'h013)) + (({mcu[375:368], 8'b0} * -24'h013)) + (({mcu[383:376], 8'b0} * -24'h02e)) + (({mcu[391:384], 8'b0} * 24'h0e7)) + (({mcu[399:392], 8'b0} * 24'h060)) + (({mcu[407:400], 8'b0} * -24'h060)) + (({mcu[415:408], 8'b0} * -24'h0e7)) + (({mcu[423:416], 8'b0} * -24'h0e7)) + (({mcu[431:424], 8'b0} * -24'h060)) + (({mcu[439:432], 8'b0} * 24'h060)) + (({mcu[447:440], 8'b0} * 24'h0e7)) + (({mcu[455:448], 8'b0} * -24'h083)) + (({mcu[463:456], 8'b0} * -24'h036)) + (({mcu[471:464], 8'b0} * 24'h036)) + (({mcu[479:472], 8'b0} * 24'h083)) + (({mcu[487:480], 8'b0} * 24'h083)) + (({mcu[495:488], 8'b0} * 24'h036)) + (({mcu[503:496], 8'b0} * -24'h036)) + (({mcu[511:504], 8'b0} * -24'h083));
	wire[47:0] cos53_term = (({mcu[7:0], 8'b0} * 24'h076)) + (({mcu[15:8], 8'b0} * -24'h01b)) + (({mcu[23:16], 8'b0} * -24'h08b)) + (({mcu[31:24], 8'b0} * -24'h04f)) + (({mcu[39:32], 8'b0} * 24'h04f)) + (({mcu[47:40], 8'b0} * 24'h08b)) + (({mcu[55:48], 8'b0} * 24'h01b)) + (({mcu[63:56], 8'b0} * -24'h076)) + (({mcu[71:64], 8'b0} * -24'h0d0)) + (({mcu[79:72], 8'b0} * 24'h030)) + (({mcu[87:80], 8'b0} * 24'h0f6)) + (({mcu[95:88], 8'b0} * 24'h08b)) + (({mcu[103:96], 8'b0} * -24'h08b)) + (({mcu[111:104], 8'b0} * -24'h0f6)) + (({mcu[119:112], 8'b0} * -24'h030)) + (({mcu[127:120], 8'b0} * 24'h0d0)) + (({mcu[135:128], 8'b0} * 24'h029)) + (({mcu[143:136], 8'b0} * -24'h009)) + (({mcu[151:144], 8'b0} * -24'h030)) + (({mcu[159:152], 8'b0} * -24'h01b)) + (({mcu[167:160], 8'b0} * 24'h01b)) + (({mcu[175:168], 8'b0} * 24'h030)) + (({mcu[183:176], 8'b0} * 24'h009)) + (({mcu[191:184], 8'b0} * -24'h029)) + (({mcu[199:192], 8'b0} * 24'h0b0)) + (({mcu[207:200], 8'b0} * -24'h029)) + (({mcu[215:208], 8'b0} * -24'h0d0)) + (({mcu[223:216], 8'b0} * -24'h076)) + (({mcu[231:224], 8'b0} * 24'h076)) + (({mcu[239:232], 8'b0} * 24'h0d0)) + (({mcu[247:240], 8'b0} * 24'h029)) + (({mcu[255:248], 8'b0} * -24'h0b0)) + (({mcu[263:256], 8'b0} * -24'h0b0)) + (({mcu[271:264], 8'b0} * 24'h029)) + (({mcu[279:272], 8'b0} * 24'h0d0)) + (({mcu[287:280], 8'b0} * 24'h076)) + (({mcu[295:288], 8'b0} * -24'h076)) + (({mcu[303:296], 8'b0} * -24'h0d0)) + (({mcu[311:304], 8'b0} * -24'h029)) + (({mcu[319:312], 8'b0} * 24'h0b0)) + (({mcu[327:320], 8'b0} * -24'h029)) + (({mcu[335:328], 8'b0} * 24'h009)) + (({mcu[343:336], 8'b0} * 24'h030)) + (({mcu[351:344], 8'b0} * 24'h01b)) + (({mcu[359:352], 8'b0} * -24'h01b)) + (({mcu[367:360], 8'b0} * -24'h030)) + (({mcu[375:368], 8'b0} * -24'h009)) + (({mcu[383:376], 8'b0} * 24'h029)) + (({mcu[391:384], 8'b0} * 24'h0d0)) + (({mcu[399:392], 8'b0} * -24'h030)) + (({mcu[407:400], 8'b0} * -24'h0f6)) + (({mcu[415:408], 8'b0} * -24'h08b)) + (({mcu[423:416], 8'b0} * 24'h08b)) + (({mcu[431:424], 8'b0} * 24'h0f6)) + (({mcu[439:432], 8'b0} * 24'h030)) + (({mcu[447:440], 8'b0} * -24'h0d0)) + (({mcu[455:448], 8'b0} * -24'h076)) + (({mcu[463:456], 8'b0} * 24'h01b)) + (({mcu[471:464], 8'b0} * 24'h08b)) + (({mcu[479:472], 8'b0} * 24'h04f)) + (({mcu[487:480], 8'b0} * -24'h04f)) + (({mcu[495:488], 8'b0} * -24'h08b)) + (({mcu[503:496], 8'b0} * -24'h01b)) + (({mcu[511:504], 8'b0} * 24'h076));
	wire[47:0] cos54_term = (({mcu[7:0], 8'b0} * 24'h064)) + (({mcu[15:8], 8'b0} * -24'h064)) + (({mcu[23:16], 8'b0} * -24'h064)) + (({mcu[31:24], 8'b0} * 24'h064)) + (({mcu[39:32], 8'b0} * 24'h064)) + (({mcu[47:40], 8'b0} * -24'h064)) + (({mcu[55:48], 8'b0} * -24'h064)) + (({mcu[63:56], 8'b0} * 24'h064)) + (({mcu[71:64], 8'b0} * -24'h0b1)) + (({mcu[79:72], 8'b0} * 24'h0b1)) + (({mcu[87:80], 8'b0} * 24'h0b1)) + (({mcu[95:88], 8'b0} * -24'h0b1)) + (({mcu[103:96], 8'b0} * -24'h0b1)) + (({mcu[111:104], 8'b0} * 24'h0b1)) + (({mcu[119:112], 8'b0} * 24'h0b1)) + (({mcu[127:120], 8'b0} * -24'h0b1)) + (({mcu[135:128], 8'b0} * 24'h023)) + (({mcu[143:136], 8'b0} * -24'h023)) + (({mcu[151:144], 8'b0} * -24'h023)) + (({mcu[159:152], 8'b0} * 24'h023)) + (({mcu[167:160], 8'b0} * 24'h023)) + (({mcu[175:168], 8'b0} * -24'h023)) + (({mcu[183:176], 8'b0} * -24'h023)) + (({mcu[191:184], 8'b0} * 24'h023)) + (({mcu[199:192], 8'b0} * 24'h096)) + (({mcu[207:200], 8'b0} * -24'h096)) + (({mcu[215:208], 8'b0} * -24'h096)) + (({mcu[223:216], 8'b0} * 24'h096)) + (({mcu[231:224], 8'b0} * 24'h096)) + (({mcu[239:232], 8'b0} * -24'h096)) + (({mcu[247:240], 8'b0} * -24'h096)) + (({mcu[255:248], 8'b0} * 24'h096)) + (({mcu[263:256], 8'b0} * -24'h096)) + (({mcu[271:264], 8'b0} * 24'h096)) + (({mcu[279:272], 8'b0} * 24'h096)) + (({mcu[287:280], 8'b0} * -24'h096)) + (({mcu[295:288], 8'b0} * -24'h096)) + (({mcu[303:296], 8'b0} * 24'h096)) + (({mcu[311:304], 8'b0} * 24'h096)) + (({mcu[319:312], 8'b0} * -24'h096)) + (({mcu[327:320], 8'b0} * -24'h023)) + (({mcu[335:328], 8'b0} * 24'h023)) + (({mcu[343:336], 8'b0} * 24'h023)) + (({mcu[351:344], 8'b0} * -24'h023)) + (({mcu[359:352], 8'b0} * -24'h023)) + (({mcu[367:360], 8'b0} * 24'h023)) + (({mcu[375:368], 8'b0} * 24'h023)) + (({mcu[383:376], 8'b0} * -24'h023)) + (({mcu[391:384], 8'b0} * 24'h0b1)) + (({mcu[399:392], 8'b0} * -24'h0b1)) + (({mcu[407:400], 8'b0} * -24'h0b1)) + (({mcu[415:408], 8'b0} * 24'h0b1)) + (({mcu[423:416], 8'b0} * 24'h0b1)) + (({mcu[431:424], 8'b0} * -24'h0b1)) + (({mcu[439:432], 8'b0} * -24'h0b1)) + (({mcu[447:440], 8'b0} * 24'h0b1)) + (({mcu[455:448], 8'b0} * -24'h064)) + (({mcu[463:456], 8'b0} * 24'h064)) + (({mcu[471:464], 8'b0} * 24'h064)) + (({mcu[479:472], 8'b0} * -24'h064)) + (({mcu[487:480], 8'b0} * -24'h064)) + (({mcu[495:488], 8'b0} * 24'h064)) + (({mcu[503:496], 8'b0} * 24'h064)) + (({mcu[511:504], 8'b0} * -24'h064));
	wire[47:0] cos55_term = (({mcu[7:0], 8'b0} * 24'h04f)) + (({mcu[15:8], 8'b0} * -24'h08b)) + (({mcu[23:16], 8'b0} * 24'h01b)) + (({mcu[31:24], 8'b0} * 24'h076)) + (({mcu[39:32], 8'b0} * -24'h076)) + (({mcu[47:40], 8'b0} * -24'h01b)) + (({mcu[55:48], 8'b0} * 24'h08b)) + (({mcu[63:56], 8'b0} * -24'h04f)) + (({mcu[71:64], 8'b0} * -24'h08b)) + (({mcu[79:72], 8'b0} * 24'h0f6)) + (({mcu[87:80], 8'b0} * -24'h030)) + (({mcu[95:88], 8'b0} * -24'h0d0)) + (({mcu[103:96], 8'b0} * 24'h0d0)) + (({mcu[111:104], 8'b0} * 24'h030)) + (({mcu[119:112], 8'b0} * -24'h0f6)) + (({mcu[127:120], 8'b0} * 24'h08b)) + (({mcu[135:128], 8'b0} * 24'h01b)) + (({mcu[143:136], 8'b0} * -24'h030)) + (({mcu[151:144], 8'b0} * 24'h009)) + (({mcu[159:152], 8'b0} * 24'h029)) + (({mcu[167:160], 8'b0} * -24'h029)) + (({mcu[175:168], 8'b0} * -24'h009)) + (({mcu[183:176], 8'b0} * 24'h030)) + (({mcu[191:184], 8'b0} * -24'h01b)) + (({mcu[199:192], 8'b0} * 24'h076)) + (({mcu[207:200], 8'b0} * -24'h0d0)) + (({mcu[215:208], 8'b0} * 24'h029)) + (({mcu[223:216], 8'b0} * 24'h0b0)) + (({mcu[231:224], 8'b0} * -24'h0b0)) + (({mcu[239:232], 8'b0} * -24'h029)) + (({mcu[247:240], 8'b0} * 24'h0d0)) + (({mcu[255:248], 8'b0} * -24'h076)) + (({mcu[263:256], 8'b0} * -24'h076)) + (({mcu[271:264], 8'b0} * 24'h0d0)) + (({mcu[279:272], 8'b0} * -24'h029)) + (({mcu[287:280], 8'b0} * -24'h0b0)) + (({mcu[295:288], 8'b0} * 24'h0b0)) + (({mcu[303:296], 8'b0} * 24'h029)) + (({mcu[311:304], 8'b0} * -24'h0d0)) + (({mcu[319:312], 8'b0} * 24'h076)) + (({mcu[327:320], 8'b0} * -24'h01b)) + (({mcu[335:328], 8'b0} * 24'h030)) + (({mcu[343:336], 8'b0} * -24'h009)) + (({mcu[351:344], 8'b0} * -24'h029)) + (({mcu[359:352], 8'b0} * 24'h029)) + (({mcu[367:360], 8'b0} * 24'h009)) + (({mcu[375:368], 8'b0} * -24'h030)) + (({mcu[383:376], 8'b0} * 24'h01b)) + (({mcu[391:384], 8'b0} * 24'h08b)) + (({mcu[399:392], 8'b0} * -24'h0f6)) + (({mcu[407:400], 8'b0} * 24'h030)) + (({mcu[415:408], 8'b0} * 24'h0d0)) + (({mcu[423:416], 8'b0} * -24'h0d0)) + (({mcu[431:424], 8'b0} * -24'h030)) + (({mcu[439:432], 8'b0} * 24'h0f6)) + (({mcu[447:440], 8'b0} * -24'h08b)) + (({mcu[455:448], 8'b0} * -24'h04f)) + (({mcu[463:456], 8'b0} * 24'h08b)) + (({mcu[471:464], 8'b0} * -24'h01b)) + (({mcu[479:472], 8'b0} * -24'h076)) + (({mcu[487:480], 8'b0} * 24'h076)) + (({mcu[495:488], 8'b0} * 24'h01b)) + (({mcu[503:496], 8'b0} * -24'h08b)) + (({mcu[511:504], 8'b0} * 24'h04f));
	wire[47:0] cos56_term = (({mcu[7:0], 8'b0} * 24'h036)) + (({mcu[15:8], 8'b0} * -24'h083)) + (({mcu[23:16], 8'b0} * 24'h083)) + (({mcu[31:24], 8'b0} * -24'h036)) + (({mcu[39:32], 8'b0} * -24'h036)) + (({mcu[47:40], 8'b0} * 24'h083)) + (({mcu[55:48], 8'b0} * -24'h083)) + (({mcu[63:56], 8'b0} * 24'h036)) + (({mcu[71:64], 8'b0} * -24'h060)) + (({mcu[79:72], 8'b0} * 24'h0e7)) + (({mcu[87:80], 8'b0} * -24'h0e7)) + (({mcu[95:88], 8'b0} * 24'h060)) + (({mcu[103:96], 8'b0} * 24'h060)) + (({mcu[111:104], 8'b0} * -24'h0e7)) + (({mcu[119:112], 8'b0} * 24'h0e7)) + (({mcu[127:120], 8'b0} * -24'h060)) + (({mcu[135:128], 8'b0} * 24'h013)) + (({mcu[143:136], 8'b0} * -24'h02e)) + (({mcu[151:144], 8'b0} * 24'h02e)) + (({mcu[159:152], 8'b0} * -24'h013)) + (({mcu[167:160], 8'b0} * -24'h013)) + (({mcu[175:168], 8'b0} * 24'h02e)) + (({mcu[183:176], 8'b0} * -24'h02e)) + (({mcu[191:184], 8'b0} * 24'h013)) + (({mcu[199:192], 8'b0} * 24'h051)) + (({mcu[207:200], 8'b0} * -24'h0c4)) + (({mcu[215:208], 8'b0} * 24'h0c4)) + (({mcu[223:216], 8'b0} * -24'h051)) + (({mcu[231:224], 8'b0} * -24'h051)) + (({mcu[239:232], 8'b0} * 24'h0c4)) + (({mcu[247:240], 8'b0} * -24'h0c4)) + (({mcu[255:248], 8'b0} * 24'h051)) + (({mcu[263:256], 8'b0} * -24'h051)) + (({mcu[271:264], 8'b0} * 24'h0c4)) + (({mcu[279:272], 8'b0} * -24'h0c4)) + (({mcu[287:280], 8'b0} * 24'h051)) + (({mcu[295:288], 8'b0} * 24'h051)) + (({mcu[303:296], 8'b0} * -24'h0c4)) + (({mcu[311:304], 8'b0} * 24'h0c4)) + (({mcu[319:312], 8'b0} * -24'h051)) + (({mcu[327:320], 8'b0} * -24'h013)) + (({mcu[335:328], 8'b0} * 24'h02e)) + (({mcu[343:336], 8'b0} * -24'h02e)) + (({mcu[351:344], 8'b0} * 24'h013)) + (({mcu[359:352], 8'b0} * 24'h013)) + (({mcu[367:360], 8'b0} * -24'h02e)) + (({mcu[375:368], 8'b0} * 24'h02e)) + (({mcu[383:376], 8'b0} * -24'h013)) + (({mcu[391:384], 8'b0} * 24'h060)) + (({mcu[399:392], 8'b0} * -24'h0e7)) + (({mcu[407:400], 8'b0} * 24'h0e7)) + (({mcu[415:408], 8'b0} * -24'h060)) + (({mcu[423:416], 8'b0} * -24'h060)) + (({mcu[431:424], 8'b0} * 24'h0e7)) + (({mcu[439:432], 8'b0} * -24'h0e7)) + (({mcu[447:440], 8'b0} * 24'h060)) + (({mcu[455:448], 8'b0} * -24'h036)) + (({mcu[463:456], 8'b0} * 24'h083)) + (({mcu[471:464], 8'b0} * -24'h083)) + (({mcu[479:472], 8'b0} * 24'h036)) + (({mcu[487:480], 8'b0} * 24'h036)) + (({mcu[495:488], 8'b0} * -24'h083)) + (({mcu[503:496], 8'b0} * 24'h083)) + (({mcu[511:504], 8'b0} * -24'h036));
	wire[47:0] cos57_term = (({mcu[7:0], 8'b0} * 24'h01b)) + (({mcu[15:8], 8'b0} * -24'h04f)) + (({mcu[23:16], 8'b0} * 24'h076)) + (({mcu[31:24], 8'b0} * -24'h08b)) + (({mcu[39:32], 8'b0} * 24'h08b)) + (({mcu[47:40], 8'b0} * -24'h076)) + (({mcu[55:48], 8'b0} * 24'h04f)) + (({mcu[63:56], 8'b0} * -24'h01b)) + (({mcu[71:64], 8'b0} * -24'h030)) + (({mcu[79:72], 8'b0} * 24'h08b)) + (({mcu[87:80], 8'b0} * -24'h0d0)) + (({mcu[95:88], 8'b0} * 24'h0f6)) + (({mcu[103:96], 8'b0} * -24'h0f6)) + (({mcu[111:104], 8'b0} * 24'h0d0)) + (({mcu[119:112], 8'b0} * -24'h08b)) + (({mcu[127:120], 8'b0} * 24'h030)) + (({mcu[135:128], 8'b0} * 24'h009)) + (({mcu[143:136], 8'b0} * -24'h01b)) + (({mcu[151:144], 8'b0} * 24'h029)) + (({mcu[159:152], 8'b0} * -24'h030)) + (({mcu[167:160], 8'b0} * 24'h030)) + (({mcu[175:168], 8'b0} * -24'h029)) + (({mcu[183:176], 8'b0} * 24'h01b)) + (({mcu[191:184], 8'b0} * -24'h009)) + (({mcu[199:192], 8'b0} * 24'h029)) + (({mcu[207:200], 8'b0} * -24'h076)) + (({mcu[215:208], 8'b0} * 24'h0b0)) + (({mcu[223:216], 8'b0} * -24'h0d0)) + (({mcu[231:224], 8'b0} * 24'h0d0)) + (({mcu[239:232], 8'b0} * -24'h0b0)) + (({mcu[247:240], 8'b0} * 24'h076)) + (({mcu[255:248], 8'b0} * -24'h029)) + (({mcu[263:256], 8'b0} * -24'h029)) + (({mcu[271:264], 8'b0} * 24'h076)) + (({mcu[279:272], 8'b0} * -24'h0b0)) + (({mcu[287:280], 8'b0} * 24'h0d0)) + (({mcu[295:288], 8'b0} * -24'h0d0)) + (({mcu[303:296], 8'b0} * 24'h0b0)) + (({mcu[311:304], 8'b0} * -24'h076)) + (({mcu[319:312], 8'b0} * 24'h029)) + (({mcu[327:320], 8'b0} * -24'h009)) + (({mcu[335:328], 8'b0} * 24'h01b)) + (({mcu[343:336], 8'b0} * -24'h029)) + (({mcu[351:344], 8'b0} * 24'h030)) + (({mcu[359:352], 8'b0} * -24'h030)) + (({mcu[367:360], 8'b0} * 24'h029)) + (({mcu[375:368], 8'b0} * -24'h01b)) + (({mcu[383:376], 8'b0} * 24'h009)) + (({mcu[391:384], 8'b0} * 24'h030)) + (({mcu[399:392], 8'b0} * -24'h08b)) + (({mcu[407:400], 8'b0} * 24'h0d0)) + (({mcu[415:408], 8'b0} * -24'h0f6)) + (({mcu[423:416], 8'b0} * 24'h0f6)) + (({mcu[431:424], 8'b0} * -24'h0d0)) + (({mcu[439:432], 8'b0} * 24'h08b)) + (({mcu[447:440], 8'b0} * -24'h030)) + (({mcu[455:448], 8'b0} * -24'h01b)) + (({mcu[463:456], 8'b0} * 24'h04f)) + (({mcu[471:464], 8'b0} * -24'h076)) + (({mcu[479:472], 8'b0} * 24'h08b)) + (({mcu[487:480], 8'b0} * -24'h08b)) + (({mcu[495:488], 8'b0} * 24'h076)) + (({mcu[503:496], 8'b0} * -24'h04f)) + (({mcu[511:504], 8'b0} * 24'h01b));
	wire[47:0] cos60_term = (({mcu[7:0], 8'b0} * 24'h062)) + (({mcu[15:8], 8'b0} * 24'h062)) + (({mcu[23:16], 8'b0} * 24'h062)) + (({mcu[31:24], 8'b0} * 24'h062)) + (({mcu[39:32], 8'b0} * 24'h062)) + (({mcu[47:40], 8'b0} * 24'h062)) + (({mcu[55:48], 8'b0} * 24'h062)) + (({mcu[63:56], 8'b0} * 24'h062)) + (({mcu[71:64], 8'b0} * -24'h0ec)) + (({mcu[79:72], 8'b0} * -24'h0ec)) + (({mcu[87:80], 8'b0} * -24'h0ec)) + (({mcu[95:88], 8'b0} * -24'h0ec)) + (({mcu[103:96], 8'b0} * -24'h0ec)) + (({mcu[111:104], 8'b0} * -24'h0ec)) + (({mcu[119:112], 8'b0} * -24'h0ec)) + (({mcu[127:120], 8'b0} * -24'h0ec)) + (({mcu[135:128], 8'b0} * 24'h0ec)) + (({mcu[143:136], 8'b0} * 24'h0ec)) + (({mcu[151:144], 8'b0} * 24'h0ec)) + (({mcu[159:152], 8'b0} * 24'h0ec)) + (({mcu[167:160], 8'b0} * 24'h0ec)) + (({mcu[175:168], 8'b0} * 24'h0ec)) + (({mcu[183:176], 8'b0} * 24'h0ec)) + (({mcu[191:184], 8'b0} * 24'h0ec)) + (({mcu[199:192], 8'b0} * -24'h062)) + (({mcu[207:200], 8'b0} * -24'h062)) + (({mcu[215:208], 8'b0} * -24'h062)) + (({mcu[223:216], 8'b0} * -24'h062)) + (({mcu[231:224], 8'b0} * -24'h062)) + (({mcu[239:232], 8'b0} * -24'h062)) + (({mcu[247:240], 8'b0} * -24'h062)) + (({mcu[255:248], 8'b0} * -24'h062)) + (({mcu[263:256], 8'b0} * -24'h062)) + (({mcu[271:264], 8'b0} * -24'h062)) + (({mcu[279:272], 8'b0} * -24'h062)) + (({mcu[287:280], 8'b0} * -24'h062)) + (({mcu[295:288], 8'b0} * -24'h062)) + (({mcu[303:296], 8'b0} * -24'h062)) + (({mcu[311:304], 8'b0} * -24'h062)) + (({mcu[319:312], 8'b0} * -24'h062)) + (({mcu[327:320], 8'b0} * 24'h0ec)) + (({mcu[335:328], 8'b0} * 24'h0ec)) + (({mcu[343:336], 8'b0} * 24'h0ec)) + (({mcu[351:344], 8'b0} * 24'h0ec)) + (({mcu[359:352], 8'b0} * 24'h0ec)) + (({mcu[367:360], 8'b0} * 24'h0ec)) + (({mcu[375:368], 8'b0} * 24'h0ec)) + (({mcu[383:376], 8'b0} * 24'h0ec)) + (({mcu[391:384], 8'b0} * -24'h0ec)) + (({mcu[399:392], 8'b0} * -24'h0ec)) + (({mcu[407:400], 8'b0} * -24'h0ec)) + (({mcu[415:408], 8'b0} * -24'h0ec)) + (({mcu[423:416], 8'b0} * -24'h0ec)) + (({mcu[431:424], 8'b0} * -24'h0ec)) + (({mcu[439:432], 8'b0} * -24'h0ec)) + (({mcu[447:440], 8'b0} * -24'h0ec)) + (({mcu[455:448], 8'b0} * 24'h062)) + (({mcu[463:456], 8'b0} * 24'h062)) + (({mcu[471:464], 8'b0} * 24'h062)) + (({mcu[479:472], 8'b0} * 24'h062)) + (({mcu[487:480], 8'b0} * 24'h062)) + (({mcu[495:488], 8'b0} * 24'h062)) + (({mcu[503:496], 8'b0} * 24'h062)) + (({mcu[511:504], 8'b0} * 24'h062));
	wire[47:0] cos61_term = (({mcu[7:0], 8'b0} * 24'h060)) + (({mcu[15:8], 8'b0} * 24'h051)) + (({mcu[23:16], 8'b0} * 24'h036)) + (({mcu[31:24], 8'b0} * 24'h013)) + (({mcu[39:32], 8'b0} * -24'h013)) + (({mcu[47:40], 8'b0} * -24'h036)) + (({mcu[55:48], 8'b0} * -24'h051)) + (({mcu[63:56], 8'b0} * -24'h060)) + (({mcu[71:64], 8'b0} * -24'h0e7)) + (({mcu[79:72], 8'b0} * -24'h0c4)) + (({mcu[87:80], 8'b0} * -24'h083)) + (({mcu[95:88], 8'b0} * -24'h02e)) + (({mcu[103:96], 8'b0} * 24'h02e)) + (({mcu[111:104], 8'b0} * 24'h083)) + (({mcu[119:112], 8'b0} * 24'h0c4)) + (({mcu[127:120], 8'b0} * 24'h0e7)) + (({mcu[135:128], 8'b0} * 24'h0e7)) + (({mcu[143:136], 8'b0} * 24'h0c4)) + (({mcu[151:144], 8'b0} * 24'h083)) + (({mcu[159:152], 8'b0} * 24'h02e)) + (({mcu[167:160], 8'b0} * -24'h02e)) + (({mcu[175:168], 8'b0} * -24'h083)) + (({mcu[183:176], 8'b0} * -24'h0c4)) + (({mcu[191:184], 8'b0} * -24'h0e7)) + (({mcu[199:192], 8'b0} * -24'h060)) + (({mcu[207:200], 8'b0} * -24'h051)) + (({mcu[215:208], 8'b0} * -24'h036)) + (({mcu[223:216], 8'b0} * -24'h013)) + (({mcu[231:224], 8'b0} * 24'h013)) + (({mcu[239:232], 8'b0} * 24'h036)) + (({mcu[247:240], 8'b0} * 24'h051)) + (({mcu[255:248], 8'b0} * 24'h060)) + (({mcu[263:256], 8'b0} * -24'h060)) + (({mcu[271:264], 8'b0} * -24'h051)) + (({mcu[279:272], 8'b0} * -24'h036)) + (({mcu[287:280], 8'b0} * -24'h013)) + (({mcu[295:288], 8'b0} * 24'h013)) + (({mcu[303:296], 8'b0} * 24'h036)) + (({mcu[311:304], 8'b0} * 24'h051)) + (({mcu[319:312], 8'b0} * 24'h060)) + (({mcu[327:320], 8'b0} * 24'h0e7)) + (({mcu[335:328], 8'b0} * 24'h0c4)) + (({mcu[343:336], 8'b0} * 24'h083)) + (({mcu[351:344], 8'b0} * 24'h02e)) + (({mcu[359:352], 8'b0} * -24'h02e)) + (({mcu[367:360], 8'b0} * -24'h083)) + (({mcu[375:368], 8'b0} * -24'h0c4)) + (({mcu[383:376], 8'b0} * -24'h0e7)) + (({mcu[391:384], 8'b0} * -24'h0e7)) + (({mcu[399:392], 8'b0} * -24'h0c4)) + (({mcu[407:400], 8'b0} * -24'h083)) + (({mcu[415:408], 8'b0} * -24'h02e)) + (({mcu[423:416], 8'b0} * 24'h02e)) + (({mcu[431:424], 8'b0} * 24'h083)) + (({mcu[439:432], 8'b0} * 24'h0c4)) + (({mcu[447:440], 8'b0} * 24'h0e7)) + (({mcu[455:448], 8'b0} * 24'h060)) + (({mcu[463:456], 8'b0} * 24'h051)) + (({mcu[471:464], 8'b0} * 24'h036)) + (({mcu[479:472], 8'b0} * 24'h013)) + (({mcu[487:480], 8'b0} * -24'h013)) + (({mcu[495:488], 8'b0} * -24'h036)) + (({mcu[503:496], 8'b0} * -24'h051)) + (({mcu[511:504], 8'b0} * -24'h060));
	wire[47:0] cos62_term = (({mcu[7:0], 8'b0} * 24'h05a)) + (({mcu[15:8], 8'b0} * 24'h025)) + (({mcu[23:16], 8'b0} * -24'h025)) + (({mcu[31:24], 8'b0} * -24'h05a)) + (({mcu[39:32], 8'b0} * -24'h05a)) + (({mcu[47:40], 8'b0} * -24'h025)) + (({mcu[55:48], 8'b0} * 24'h025)) + (({mcu[63:56], 8'b0} * 24'h05a)) + (({mcu[71:64], 8'b0} * -24'h0da)) + (({mcu[79:72], 8'b0} * -24'h05a)) + (({mcu[87:80], 8'b0} * 24'h05a)) + (({mcu[95:88], 8'b0} * 24'h0da)) + (({mcu[103:96], 8'b0} * 24'h0da)) + (({mcu[111:104], 8'b0} * 24'h05a)) + (({mcu[119:112], 8'b0} * -24'h05a)) + (({mcu[127:120], 8'b0} * -24'h0da)) + (({mcu[135:128], 8'b0} * 24'h0da)) + (({mcu[143:136], 8'b0} * 24'h05a)) + (({mcu[151:144], 8'b0} * -24'h05a)) + (({mcu[159:152], 8'b0} * -24'h0da)) + (({mcu[167:160], 8'b0} * -24'h0da)) + (({mcu[175:168], 8'b0} * -24'h05a)) + (({mcu[183:176], 8'b0} * 24'h05a)) + (({mcu[191:184], 8'b0} * 24'h0da)) + (({mcu[199:192], 8'b0} * -24'h05a)) + (({mcu[207:200], 8'b0} * -24'h025)) + (({mcu[215:208], 8'b0} * 24'h025)) + (({mcu[223:216], 8'b0} * 24'h05a)) + (({mcu[231:224], 8'b0} * 24'h05a)) + (({mcu[239:232], 8'b0} * 24'h025)) + (({mcu[247:240], 8'b0} * -24'h025)) + (({mcu[255:248], 8'b0} * -24'h05a)) + (({mcu[263:256], 8'b0} * -24'h05a)) + (({mcu[271:264], 8'b0} * -24'h025)) + (({mcu[279:272], 8'b0} * 24'h025)) + (({mcu[287:280], 8'b0} * 24'h05a)) + (({mcu[295:288], 8'b0} * 24'h05a)) + (({mcu[303:296], 8'b0} * 24'h025)) + (({mcu[311:304], 8'b0} * -24'h025)) + (({mcu[319:312], 8'b0} * -24'h05a)) + (({mcu[327:320], 8'b0} * 24'h0da)) + (({mcu[335:328], 8'b0} * 24'h05a)) + (({mcu[343:336], 8'b0} * -24'h05a)) + (({mcu[351:344], 8'b0} * -24'h0da)) + (({mcu[359:352], 8'b0} * -24'h0da)) + (({mcu[367:360], 8'b0} * -24'h05a)) + (({mcu[375:368], 8'b0} * 24'h05a)) + (({mcu[383:376], 8'b0} * 24'h0da)) + (({mcu[391:384], 8'b0} * -24'h0da)) + (({mcu[399:392], 8'b0} * -24'h05a)) + (({mcu[407:400], 8'b0} * 24'h05a)) + (({mcu[415:408], 8'b0} * 24'h0da)) + (({mcu[423:416], 8'b0} * 24'h0da)) + (({mcu[431:424], 8'b0} * 24'h05a)) + (({mcu[439:432], 8'b0} * -24'h05a)) + (({mcu[447:440], 8'b0} * -24'h0da)) + (({mcu[455:448], 8'b0} * 24'h05a)) + (({mcu[463:456], 8'b0} * 24'h025)) + (({mcu[471:464], 8'b0} * -24'h025)) + (({mcu[479:472], 8'b0} * -24'h05a)) + (({mcu[487:480], 8'b0} * -24'h05a)) + (({mcu[495:488], 8'b0} * -24'h025)) + (({mcu[503:496], 8'b0} * 24'h025)) + (({mcu[511:504], 8'b0} * 24'h05a));
	wire[47:0] cos63_term = (({mcu[7:0], 8'b0} * 24'h051)) + (({mcu[15:8], 8'b0} * -24'h013)) + (({mcu[23:16], 8'b0} * -24'h060)) + (({mcu[31:24], 8'b0} * -24'h036)) + (({mcu[39:32], 8'b0} * 24'h036)) + (({mcu[47:40], 8'b0} * 24'h060)) + (({mcu[55:48], 8'b0} * 24'h013)) + (({mcu[63:56], 8'b0} * -24'h051)) + (({mcu[71:64], 8'b0} * -24'h0c4)) + (({mcu[79:72], 8'b0} * 24'h02e)) + (({mcu[87:80], 8'b0} * 24'h0e7)) + (({mcu[95:88], 8'b0} * 24'h083)) + (({mcu[103:96], 8'b0} * -24'h083)) + (({mcu[111:104], 8'b0} * -24'h0e7)) + (({mcu[119:112], 8'b0} * -24'h02e)) + (({mcu[127:120], 8'b0} * 24'h0c4)) + (({mcu[135:128], 8'b0} * 24'h0c4)) + (({mcu[143:136], 8'b0} * -24'h02e)) + (({mcu[151:144], 8'b0} * -24'h0e7)) + (({mcu[159:152], 8'b0} * -24'h083)) + (({mcu[167:160], 8'b0} * 24'h083)) + (({mcu[175:168], 8'b0} * 24'h0e7)) + (({mcu[183:176], 8'b0} * 24'h02e)) + (({mcu[191:184], 8'b0} * -24'h0c4)) + (({mcu[199:192], 8'b0} * -24'h051)) + (({mcu[207:200], 8'b0} * 24'h013)) + (({mcu[215:208], 8'b0} * 24'h060)) + (({mcu[223:216], 8'b0} * 24'h036)) + (({mcu[231:224], 8'b0} * -24'h036)) + (({mcu[239:232], 8'b0} * -24'h060)) + (({mcu[247:240], 8'b0} * -24'h013)) + (({mcu[255:248], 8'b0} * 24'h051)) + (({mcu[263:256], 8'b0} * -24'h051)) + (({mcu[271:264], 8'b0} * 24'h013)) + (({mcu[279:272], 8'b0} * 24'h060)) + (({mcu[287:280], 8'b0} * 24'h036)) + (({mcu[295:288], 8'b0} * -24'h036)) + (({mcu[303:296], 8'b0} * -24'h060)) + (({mcu[311:304], 8'b0} * -24'h013)) + (({mcu[319:312], 8'b0} * 24'h051)) + (({mcu[327:320], 8'b0} * 24'h0c4)) + (({mcu[335:328], 8'b0} * -24'h02e)) + (({mcu[343:336], 8'b0} * -24'h0e7)) + (({mcu[351:344], 8'b0} * -24'h083)) + (({mcu[359:352], 8'b0} * 24'h083)) + (({mcu[367:360], 8'b0} * 24'h0e7)) + (({mcu[375:368], 8'b0} * 24'h02e)) + (({mcu[383:376], 8'b0} * -24'h0c4)) + (({mcu[391:384], 8'b0} * -24'h0c4)) + (({mcu[399:392], 8'b0} * 24'h02e)) + (({mcu[407:400], 8'b0} * 24'h0e7)) + (({mcu[415:408], 8'b0} * 24'h083)) + (({mcu[423:416], 8'b0} * -24'h083)) + (({mcu[431:424], 8'b0} * -24'h0e7)) + (({mcu[439:432], 8'b0} * -24'h02e)) + (({mcu[447:440], 8'b0} * 24'h0c4)) + (({mcu[455:448], 8'b0} * 24'h051)) + (({mcu[463:456], 8'b0} * -24'h013)) + (({mcu[471:464], 8'b0} * -24'h060)) + (({mcu[479:472], 8'b0} * -24'h036)) + (({mcu[487:480], 8'b0} * 24'h036)) + (({mcu[495:488], 8'b0} * 24'h060)) + (({mcu[503:496], 8'b0} * 24'h013)) + (({mcu[511:504], 8'b0} * -24'h051));
	wire[47:0] cos64_term = (({mcu[7:0], 8'b0} * 24'h045)) + (({mcu[15:8], 8'b0} * -24'h045)) + (({mcu[23:16], 8'b0} * -24'h045)) + (({mcu[31:24], 8'b0} * 24'h045)) + (({mcu[39:32], 8'b0} * 24'h045)) + (({mcu[47:40], 8'b0} * -24'h045)) + (({mcu[55:48], 8'b0} * -24'h045)) + (({mcu[63:56], 8'b0} * 24'h045)) + (({mcu[71:64], 8'b0} * -24'h0a7)) + (({mcu[79:72], 8'b0} * 24'h0a7)) + (({mcu[87:80], 8'b0} * 24'h0a7)) + (({mcu[95:88], 8'b0} * -24'h0a7)) + (({mcu[103:96], 8'b0} * -24'h0a7)) + (({mcu[111:104], 8'b0} * 24'h0a7)) + (({mcu[119:112], 8'b0} * 24'h0a7)) + (({mcu[127:120], 8'b0} * -24'h0a7)) + (({mcu[135:128], 8'b0} * 24'h0a7)) + (({mcu[143:136], 8'b0} * -24'h0a7)) + (({mcu[151:144], 8'b0} * -24'h0a7)) + (({mcu[159:152], 8'b0} * 24'h0a7)) + (({mcu[167:160], 8'b0} * 24'h0a7)) + (({mcu[175:168], 8'b0} * -24'h0a7)) + (({mcu[183:176], 8'b0} * -24'h0a7)) + (({mcu[191:184], 8'b0} * 24'h0a7)) + (({mcu[199:192], 8'b0} * -24'h045)) + (({mcu[207:200], 8'b0} * 24'h045)) + (({mcu[215:208], 8'b0} * 24'h045)) + (({mcu[223:216], 8'b0} * -24'h045)) + (({mcu[231:224], 8'b0} * -24'h045)) + (({mcu[239:232], 8'b0} * 24'h045)) + (({mcu[247:240], 8'b0} * 24'h045)) + (({mcu[255:248], 8'b0} * -24'h045)) + (({mcu[263:256], 8'b0} * -24'h045)) + (({mcu[271:264], 8'b0} * 24'h045)) + (({mcu[279:272], 8'b0} * 24'h045)) + (({mcu[287:280], 8'b0} * -24'h045)) + (({mcu[295:288], 8'b0} * -24'h045)) + (({mcu[303:296], 8'b0} * 24'h045)) + (({mcu[311:304], 8'b0} * 24'h045)) + (({mcu[319:312], 8'b0} * -24'h045)) + (({mcu[327:320], 8'b0} * 24'h0a7)) + (({mcu[335:328], 8'b0} * -24'h0a7)) + (({mcu[343:336], 8'b0} * -24'h0a7)) + (({mcu[351:344], 8'b0} * 24'h0a7)) + (({mcu[359:352], 8'b0} * 24'h0a7)) + (({mcu[367:360], 8'b0} * -24'h0a7)) + (({mcu[375:368], 8'b0} * -24'h0a7)) + (({mcu[383:376], 8'b0} * 24'h0a7)) + (({mcu[391:384], 8'b0} * -24'h0a7)) + (({mcu[399:392], 8'b0} * 24'h0a7)) + (({mcu[407:400], 8'b0} * 24'h0a7)) + (({mcu[415:408], 8'b0} * -24'h0a7)) + (({mcu[423:416], 8'b0} * -24'h0a7)) + (({mcu[431:424], 8'b0} * 24'h0a7)) + (({mcu[439:432], 8'b0} * 24'h0a7)) + (({mcu[447:440], 8'b0} * -24'h0a7)) + (({mcu[455:448], 8'b0} * 24'h045)) + (({mcu[463:456], 8'b0} * -24'h045)) + (({mcu[471:464], 8'b0} * -24'h045)) + (({mcu[479:472], 8'b0} * 24'h045)) + (({mcu[487:480], 8'b0} * 24'h045)) + (({mcu[495:488], 8'b0} * -24'h045)) + (({mcu[503:496], 8'b0} * -24'h045)) + (({mcu[511:504], 8'b0} * 24'h045));
	wire[47:0] cos65_term = (({mcu[7:0], 8'b0} * 24'h036)) + (({mcu[15:8], 8'b0} * -24'h060)) + (({mcu[23:16], 8'b0} * 24'h013)) + (({mcu[31:24], 8'b0} * 24'h051)) + (({mcu[39:32], 8'b0} * -24'h051)) + (({mcu[47:40], 8'b0} * -24'h013)) + (({mcu[55:48], 8'b0} * 24'h060)) + (({mcu[63:56], 8'b0} * -24'h036)) + (({mcu[71:64], 8'b0} * -24'h083)) + (({mcu[79:72], 8'b0} * 24'h0e7)) + (({mcu[87:80], 8'b0} * -24'h02e)) + (({mcu[95:88], 8'b0} * -24'h0c4)) + (({mcu[103:96], 8'b0} * 24'h0c4)) + (({mcu[111:104], 8'b0} * 24'h02e)) + (({mcu[119:112], 8'b0} * -24'h0e7)) + (({mcu[127:120], 8'b0} * 24'h083)) + (({mcu[135:128], 8'b0} * 24'h083)) + (({mcu[143:136], 8'b0} * -24'h0e7)) + (({mcu[151:144], 8'b0} * 24'h02e)) + (({mcu[159:152], 8'b0} * 24'h0c4)) + (({mcu[167:160], 8'b0} * -24'h0c4)) + (({mcu[175:168], 8'b0} * -24'h02e)) + (({mcu[183:176], 8'b0} * 24'h0e7)) + (({mcu[191:184], 8'b0} * -24'h083)) + (({mcu[199:192], 8'b0} * -24'h036)) + (({mcu[207:200], 8'b0} * 24'h060)) + (({mcu[215:208], 8'b0} * -24'h013)) + (({mcu[223:216], 8'b0} * -24'h051)) + (({mcu[231:224], 8'b0} * 24'h051)) + (({mcu[239:232], 8'b0} * 24'h013)) + (({mcu[247:240], 8'b0} * -24'h060)) + (({mcu[255:248], 8'b0} * 24'h036)) + (({mcu[263:256], 8'b0} * -24'h036)) + (({mcu[271:264], 8'b0} * 24'h060)) + (({mcu[279:272], 8'b0} * -24'h013)) + (({mcu[287:280], 8'b0} * -24'h051)) + (({mcu[295:288], 8'b0} * 24'h051)) + (({mcu[303:296], 8'b0} * 24'h013)) + (({mcu[311:304], 8'b0} * -24'h060)) + (({mcu[319:312], 8'b0} * 24'h036)) + (({mcu[327:320], 8'b0} * 24'h083)) + (({mcu[335:328], 8'b0} * -24'h0e7)) + (({mcu[343:336], 8'b0} * 24'h02e)) + (({mcu[351:344], 8'b0} * 24'h0c4)) + (({mcu[359:352], 8'b0} * -24'h0c4)) + (({mcu[367:360], 8'b0} * -24'h02e)) + (({mcu[375:368], 8'b0} * 24'h0e7)) + (({mcu[383:376], 8'b0} * -24'h083)) + (({mcu[391:384], 8'b0} * -24'h083)) + (({mcu[399:392], 8'b0} * 24'h0e7)) + (({mcu[407:400], 8'b0} * -24'h02e)) + (({mcu[415:408], 8'b0} * -24'h0c4)) + (({mcu[423:416], 8'b0} * 24'h0c4)) + (({mcu[431:424], 8'b0} * 24'h02e)) + (({mcu[439:432], 8'b0} * -24'h0e7)) + (({mcu[447:440], 8'b0} * 24'h083)) + (({mcu[455:448], 8'b0} * 24'h036)) + (({mcu[463:456], 8'b0} * -24'h060)) + (({mcu[471:464], 8'b0} * 24'h013)) + (({mcu[479:472], 8'b0} * 24'h051)) + (({mcu[487:480], 8'b0} * -24'h051)) + (({mcu[495:488], 8'b0} * -24'h013)) + (({mcu[503:496], 8'b0} * 24'h060)) + (({mcu[511:504], 8'b0} * -24'h036));
	wire[47:0] cos66_term = (({mcu[7:0], 8'b0} * 24'h025)) + (({mcu[15:8], 8'b0} * -24'h05a)) + (({mcu[23:16], 8'b0} * 24'h05a)) + (({mcu[31:24], 8'b0} * -24'h025)) + (({mcu[39:32], 8'b0} * -24'h025)) + (({mcu[47:40], 8'b0} * 24'h05a)) + (({mcu[55:48], 8'b0} * -24'h05a)) + (({mcu[63:56], 8'b0} * 24'h025)) + (({mcu[71:64], 8'b0} * -24'h05a)) + (({mcu[79:72], 8'b0} * 24'h0da)) + (({mcu[87:80], 8'b0} * -24'h0da)) + (({mcu[95:88], 8'b0} * 24'h05a)) + (({mcu[103:96], 8'b0} * 24'h05a)) + (({mcu[111:104], 8'b0} * -24'h0da)) + (({mcu[119:112], 8'b0} * 24'h0da)) + (({mcu[127:120], 8'b0} * -24'h05a)) + (({mcu[135:128], 8'b0} * 24'h05a)) + (({mcu[143:136], 8'b0} * -24'h0da)) + (({mcu[151:144], 8'b0} * 24'h0da)) + (({mcu[159:152], 8'b0} * -24'h05a)) + (({mcu[167:160], 8'b0} * -24'h05a)) + (({mcu[175:168], 8'b0} * 24'h0da)) + (({mcu[183:176], 8'b0} * -24'h0da)) + (({mcu[191:184], 8'b0} * 24'h05a)) + (({mcu[199:192], 8'b0} * -24'h025)) + (({mcu[207:200], 8'b0} * 24'h05a)) + (({mcu[215:208], 8'b0} * -24'h05a)) + (({mcu[223:216], 8'b0} * 24'h025)) + (({mcu[231:224], 8'b0} * 24'h025)) + (({mcu[239:232], 8'b0} * -24'h05a)) + (({mcu[247:240], 8'b0} * 24'h05a)) + (({mcu[255:248], 8'b0} * -24'h025)) + (({mcu[263:256], 8'b0} * -24'h025)) + (({mcu[271:264], 8'b0} * 24'h05a)) + (({mcu[279:272], 8'b0} * -24'h05a)) + (({mcu[287:280], 8'b0} * 24'h025)) + (({mcu[295:288], 8'b0} * 24'h025)) + (({mcu[303:296], 8'b0} * -24'h05a)) + (({mcu[311:304], 8'b0} * 24'h05a)) + (({mcu[319:312], 8'b0} * -24'h025)) + (({mcu[327:320], 8'b0} * 24'h05a)) + (({mcu[335:328], 8'b0} * -24'h0da)) + (({mcu[343:336], 8'b0} * 24'h0da)) + (({mcu[351:344], 8'b0} * -24'h05a)) + (({mcu[359:352], 8'b0} * -24'h05a)) + (({mcu[367:360], 8'b0} * 24'h0da)) + (({mcu[375:368], 8'b0} * -24'h0da)) + (({mcu[383:376], 8'b0} * 24'h05a)) + (({mcu[391:384], 8'b0} * -24'h05a)) + (({mcu[399:392], 8'b0} * 24'h0da)) + (({mcu[407:400], 8'b0} * -24'h0da)) + (({mcu[415:408], 8'b0} * 24'h05a)) + (({mcu[423:416], 8'b0} * 24'h05a)) + (({mcu[431:424], 8'b0} * -24'h0da)) + (({mcu[439:432], 8'b0} * 24'h0da)) + (({mcu[447:440], 8'b0} * -24'h05a)) + (({mcu[455:448], 8'b0} * 24'h025)) + (({mcu[463:456], 8'b0} * -24'h05a)) + (({mcu[471:464], 8'b0} * 24'h05a)) + (({mcu[479:472], 8'b0} * -24'h025)) + (({mcu[487:480], 8'b0} * -24'h025)) + (({mcu[495:488], 8'b0} * 24'h05a)) + (({mcu[503:496], 8'b0} * -24'h05a)) + (({mcu[511:504], 8'b0} * 24'h025));
	wire[47:0] cos67_term = (({mcu[7:0], 8'b0} * 24'h013)) + (({mcu[15:8], 8'b0} * -24'h036)) + (({mcu[23:16], 8'b0} * 24'h051)) + (({mcu[31:24], 8'b0} * -24'h060)) + (({mcu[39:32], 8'b0} * 24'h060)) + (({mcu[47:40], 8'b0} * -24'h051)) + (({mcu[55:48], 8'b0} * 24'h036)) + (({mcu[63:56], 8'b0} * -24'h013)) + (({mcu[71:64], 8'b0} * -24'h02e)) + (({mcu[79:72], 8'b0} * 24'h083)) + (({mcu[87:80], 8'b0} * -24'h0c4)) + (({mcu[95:88], 8'b0} * 24'h0e7)) + (({mcu[103:96], 8'b0} * -24'h0e7)) + (({mcu[111:104], 8'b0} * 24'h0c4)) + (({mcu[119:112], 8'b0} * -24'h083)) + (({mcu[127:120], 8'b0} * 24'h02e)) + (({mcu[135:128], 8'b0} * 24'h02e)) + (({mcu[143:136], 8'b0} * -24'h083)) + (({mcu[151:144], 8'b0} * 24'h0c4)) + (({mcu[159:152], 8'b0} * -24'h0e7)) + (({mcu[167:160], 8'b0} * 24'h0e7)) + (({mcu[175:168], 8'b0} * -24'h0c4)) + (({mcu[183:176], 8'b0} * 24'h083)) + (({mcu[191:184], 8'b0} * -24'h02e)) + (({mcu[199:192], 8'b0} * -24'h013)) + (({mcu[207:200], 8'b0} * 24'h036)) + (({mcu[215:208], 8'b0} * -24'h051)) + (({mcu[223:216], 8'b0} * 24'h060)) + (({mcu[231:224], 8'b0} * -24'h060)) + (({mcu[239:232], 8'b0} * 24'h051)) + (({mcu[247:240], 8'b0} * -24'h036)) + (({mcu[255:248], 8'b0} * 24'h013)) + (({mcu[263:256], 8'b0} * -24'h013)) + (({mcu[271:264], 8'b0} * 24'h036)) + (({mcu[279:272], 8'b0} * -24'h051)) + (({mcu[287:280], 8'b0} * 24'h060)) + (({mcu[295:288], 8'b0} * -24'h060)) + (({mcu[303:296], 8'b0} * 24'h051)) + (({mcu[311:304], 8'b0} * -24'h036)) + (({mcu[319:312], 8'b0} * 24'h013)) + (({mcu[327:320], 8'b0} * 24'h02e)) + (({mcu[335:328], 8'b0} * -24'h083)) + (({mcu[343:336], 8'b0} * 24'h0c4)) + (({mcu[351:344], 8'b0} * -24'h0e7)) + (({mcu[359:352], 8'b0} * 24'h0e7)) + (({mcu[367:360], 8'b0} * -24'h0c4)) + (({mcu[375:368], 8'b0} * 24'h083)) + (({mcu[383:376], 8'b0} * -24'h02e)) + (({mcu[391:384], 8'b0} * -24'h02e)) + (({mcu[399:392], 8'b0} * 24'h083)) + (({mcu[407:400], 8'b0} * -24'h0c4)) + (({mcu[415:408], 8'b0} * 24'h0e7)) + (({mcu[423:416], 8'b0} * -24'h0e7)) + (({mcu[431:424], 8'b0} * 24'h0c4)) + (({mcu[439:432], 8'b0} * -24'h083)) + (({mcu[447:440], 8'b0} * 24'h02e)) + (({mcu[455:448], 8'b0} * 24'h013)) + (({mcu[463:456], 8'b0} * -24'h036)) + (({mcu[471:464], 8'b0} * 24'h051)) + (({mcu[479:472], 8'b0} * -24'h060)) + (({mcu[487:480], 8'b0} * 24'h060)) + (({mcu[495:488], 8'b0} * -24'h051)) + (({mcu[503:496], 8'b0} * 24'h036)) + (({mcu[511:504], 8'b0} * -24'h013));
	wire[47:0] cos70_term = (({mcu[7:0], 8'b0} * 24'h031)) + (({mcu[15:8], 8'b0} * 24'h031)) + (({mcu[23:16], 8'b0} * 24'h031)) + (({mcu[31:24], 8'b0} * 24'h031)) + (({mcu[39:32], 8'b0} * 24'h031)) + (({mcu[47:40], 8'b0} * 24'h031)) + (({mcu[55:48], 8'b0} * 24'h031)) + (({mcu[63:56], 8'b0} * 24'h031)) + (({mcu[71:64], 8'b0} * -24'h08e)) + (({mcu[79:72], 8'b0} * -24'h08e)) + (({mcu[87:80], 8'b0} * -24'h08e)) + (({mcu[95:88], 8'b0} * -24'h08e)) + (({mcu[103:96], 8'b0} * -24'h08e)) + (({mcu[111:104], 8'b0} * -24'h08e)) + (({mcu[119:112], 8'b0} * -24'h08e)) + (({mcu[127:120], 8'b0} * -24'h08e)) + (({mcu[135:128], 8'b0} * 24'h0d4)) + (({mcu[143:136], 8'b0} * 24'h0d4)) + (({mcu[151:144], 8'b0} * 24'h0d4)) + (({mcu[159:152], 8'b0} * 24'h0d4)) + (({mcu[167:160], 8'b0} * 24'h0d4)) + (({mcu[175:168], 8'b0} * 24'h0d4)) + (({mcu[183:176], 8'b0} * 24'h0d4)) + (({mcu[191:184], 8'b0} * 24'h0d4)) + (({mcu[199:192], 8'b0} * -24'h0fb)) + (({mcu[207:200], 8'b0} * -24'h0fb)) + (({mcu[215:208], 8'b0} * -24'h0fb)) + (({mcu[223:216], 8'b0} * -24'h0fb)) + (({mcu[231:224], 8'b0} * -24'h0fb)) + (({mcu[239:232], 8'b0} * -24'h0fb)) + (({mcu[247:240], 8'b0} * -24'h0fb)) + (({mcu[255:248], 8'b0} * -24'h0fb)) + (({mcu[263:256], 8'b0} * 24'h0fb)) + (({mcu[271:264], 8'b0} * 24'h0fb)) + (({mcu[279:272], 8'b0} * 24'h0fb)) + (({mcu[287:280], 8'b0} * 24'h0fb)) + (({mcu[295:288], 8'b0} * 24'h0fb)) + (({mcu[303:296], 8'b0} * 24'h0fb)) + (({mcu[311:304], 8'b0} * 24'h0fb)) + (({mcu[319:312], 8'b0} * 24'h0fb)) + (({mcu[327:320], 8'b0} * -24'h0d4)) + (({mcu[335:328], 8'b0} * -24'h0d4)) + (({mcu[343:336], 8'b0} * -24'h0d4)) + (({mcu[351:344], 8'b0} * -24'h0d4)) + (({mcu[359:352], 8'b0} * -24'h0d4)) + (({mcu[367:360], 8'b0} * -24'h0d4)) + (({mcu[375:368], 8'b0} * -24'h0d4)) + (({mcu[383:376], 8'b0} * -24'h0d4)) + (({mcu[391:384], 8'b0} * 24'h08e)) + (({mcu[399:392], 8'b0} * 24'h08e)) + (({mcu[407:400], 8'b0} * 24'h08e)) + (({mcu[415:408], 8'b0} * 24'h08e)) + (({mcu[423:416], 8'b0} * 24'h08e)) + (({mcu[431:424], 8'b0} * 24'h08e)) + (({mcu[439:432], 8'b0} * 24'h08e)) + (({mcu[447:440], 8'b0} * 24'h08e)) + (({mcu[455:448], 8'b0} * -24'h031)) + (({mcu[463:456], 8'b0} * -24'h031)) + (({mcu[471:464], 8'b0} * -24'h031)) + (({mcu[479:472], 8'b0} * -24'h031)) + (({mcu[487:480], 8'b0} * -24'h031)) + (({mcu[495:488], 8'b0} * -24'h031)) + (({mcu[503:496], 8'b0} * -24'h031)) + (({mcu[511:504], 8'b0} * -24'h031));
	wire[47:0] cos71_term = (({mcu[7:0], 8'b0} * 24'h030)) + (({mcu[15:8], 8'b0} * 24'h029)) + (({mcu[23:16], 8'b0} * 24'h01b)) + (({mcu[31:24], 8'b0} * 24'h009)) + (({mcu[39:32], 8'b0} * -24'h009)) + (({mcu[47:40], 8'b0} * -24'h01b)) + (({mcu[55:48], 8'b0} * -24'h029)) + (({mcu[63:56], 8'b0} * -24'h030)) + (({mcu[71:64], 8'b0} * -24'h08b)) + (({mcu[79:72], 8'b0} * -24'h076)) + (({mcu[87:80], 8'b0} * -24'h04f)) + (({mcu[95:88], 8'b0} * -24'h01b)) + (({mcu[103:96], 8'b0} * 24'h01b)) + (({mcu[111:104], 8'b0} * 24'h04f)) + (({mcu[119:112], 8'b0} * 24'h076)) + (({mcu[127:120], 8'b0} * 24'h08b)) + (({mcu[135:128], 8'b0} * 24'h0d0)) + (({mcu[143:136], 8'b0} * 24'h0b0)) + (({mcu[151:144], 8'b0} * 24'h076)) + (({mcu[159:152], 8'b0} * 24'h029)) + (({mcu[167:160], 8'b0} * -24'h029)) + (({mcu[175:168], 8'b0} * -24'h076)) + (({mcu[183:176], 8'b0} * -24'h0b0)) + (({mcu[191:184], 8'b0} * -24'h0d0)) + (({mcu[199:192], 8'b0} * -24'h0f6)) + (({mcu[207:200], 8'b0} * -24'h0d0)) + (({mcu[215:208], 8'b0} * -24'h08b)) + (({mcu[223:216], 8'b0} * -24'h030)) + (({mcu[231:224], 8'b0} * 24'h030)) + (({mcu[239:232], 8'b0} * 24'h08b)) + (({mcu[247:240], 8'b0} * 24'h0d0)) + (({mcu[255:248], 8'b0} * 24'h0f6)) + (({mcu[263:256], 8'b0} * 24'h0f6)) + (({mcu[271:264], 8'b0} * 24'h0d0)) + (({mcu[279:272], 8'b0} * 24'h08b)) + (({mcu[287:280], 8'b0} * 24'h030)) + (({mcu[295:288], 8'b0} * -24'h030)) + (({mcu[303:296], 8'b0} * -24'h08b)) + (({mcu[311:304], 8'b0} * -24'h0d0)) + (({mcu[319:312], 8'b0} * -24'h0f6)) + (({mcu[327:320], 8'b0} * -24'h0d0)) + (({mcu[335:328], 8'b0} * -24'h0b0)) + (({mcu[343:336], 8'b0} * -24'h076)) + (({mcu[351:344], 8'b0} * -24'h029)) + (({mcu[359:352], 8'b0} * 24'h029)) + (({mcu[367:360], 8'b0} * 24'h076)) + (({mcu[375:368], 8'b0} * 24'h0b0)) + (({mcu[383:376], 8'b0} * 24'h0d0)) + (({mcu[391:384], 8'b0} * 24'h08b)) + (({mcu[399:392], 8'b0} * 24'h076)) + (({mcu[407:400], 8'b0} * 24'h04f)) + (({mcu[415:408], 8'b0} * 24'h01b)) + (({mcu[423:416], 8'b0} * -24'h01b)) + (({mcu[431:424], 8'b0} * -24'h04f)) + (({mcu[439:432], 8'b0} * -24'h076)) + (({mcu[447:440], 8'b0} * -24'h08b)) + (({mcu[455:448], 8'b0} * -24'h030)) + (({mcu[463:456], 8'b0} * -24'h029)) + (({mcu[471:464], 8'b0} * -24'h01b)) + (({mcu[479:472], 8'b0} * -24'h009)) + (({mcu[487:480], 8'b0} * 24'h009)) + (({mcu[495:488], 8'b0} * 24'h01b)) + (({mcu[503:496], 8'b0} * 24'h029)) + (({mcu[511:504], 8'b0} * 24'h030));
	wire[47:0] cos72_term = (({mcu[7:0], 8'b0} * 24'h02e)) + (({mcu[15:8], 8'b0} * 24'h013)) + (({mcu[23:16], 8'b0} * -24'h013)) + (({mcu[31:24], 8'b0} * -24'h02e)) + (({mcu[39:32], 8'b0} * -24'h02e)) + (({mcu[47:40], 8'b0} * -24'h013)) + (({mcu[55:48], 8'b0} * 24'h013)) + (({mcu[63:56], 8'b0} * 24'h02e)) + (({mcu[71:64], 8'b0} * -24'h083)) + (({mcu[79:72], 8'b0} * -24'h036)) + (({mcu[87:80], 8'b0} * 24'h036)) + (({mcu[95:88], 8'b0} * 24'h083)) + (({mcu[103:96], 8'b0} * 24'h083)) + (({mcu[111:104], 8'b0} * 24'h036)) + (({mcu[119:112], 8'b0} * -24'h036)) + (({mcu[127:120], 8'b0} * -24'h083)) + (({mcu[135:128], 8'b0} * 24'h0c4)) + (({mcu[143:136], 8'b0} * 24'h051)) + (({mcu[151:144], 8'b0} * -24'h051)) + (({mcu[159:152], 8'b0} * -24'h0c4)) + (({mcu[167:160], 8'b0} * -24'h0c4)) + (({mcu[175:168], 8'b0} * -24'h051)) + (({mcu[183:176], 8'b0} * 24'h051)) + (({mcu[191:184], 8'b0} * 24'h0c4)) + (({mcu[199:192], 8'b0} * -24'h0e7)) + (({mcu[207:200], 8'b0} * -24'h060)) + (({mcu[215:208], 8'b0} * 24'h060)) + (({mcu[223:216], 8'b0} * 24'h0e7)) + (({mcu[231:224], 8'b0} * 24'h0e7)) + (({mcu[239:232], 8'b0} * 24'h060)) + (({mcu[247:240], 8'b0} * -24'h060)) + (({mcu[255:248], 8'b0} * -24'h0e7)) + (({mcu[263:256], 8'b0} * 24'h0e7)) + (({mcu[271:264], 8'b0} * 24'h060)) + (({mcu[279:272], 8'b0} * -24'h060)) + (({mcu[287:280], 8'b0} * -24'h0e7)) + (({mcu[295:288], 8'b0} * -24'h0e7)) + (({mcu[303:296], 8'b0} * -24'h060)) + (({mcu[311:304], 8'b0} * 24'h060)) + (({mcu[319:312], 8'b0} * 24'h0e7)) + (({mcu[327:320], 8'b0} * -24'h0c4)) + (({mcu[335:328], 8'b0} * -24'h051)) + (({mcu[343:336], 8'b0} * 24'h051)) + (({mcu[351:344], 8'b0} * 24'h0c4)) + (({mcu[359:352], 8'b0} * 24'h0c4)) + (({mcu[367:360], 8'b0} * 24'h051)) + (({mcu[375:368], 8'b0} * -24'h051)) + (({mcu[383:376], 8'b0} * -24'h0c4)) + (({mcu[391:384], 8'b0} * 24'h083)) + (({mcu[399:392], 8'b0} * 24'h036)) + (({mcu[407:400], 8'b0} * -24'h036)) + (({mcu[415:408], 8'b0} * -24'h083)) + (({mcu[423:416], 8'b0} * -24'h083)) + (({mcu[431:424], 8'b0} * -24'h036)) + (({mcu[439:432], 8'b0} * 24'h036)) + (({mcu[447:440], 8'b0} * 24'h083)) + (({mcu[455:448], 8'b0} * -24'h02e)) + (({mcu[463:456], 8'b0} * -24'h013)) + (({mcu[471:464], 8'b0} * 24'h013)) + (({mcu[479:472], 8'b0} * 24'h02e)) + (({mcu[487:480], 8'b0} * 24'h02e)) + (({mcu[495:488], 8'b0} * 24'h013)) + (({mcu[503:496], 8'b0} * -24'h013)) + (({mcu[511:504], 8'b0} * -24'h02e));
	wire[47:0] cos73_term = (({mcu[7:0], 8'b0} * 24'h029)) + (({mcu[15:8], 8'b0} * -24'h009)) + (({mcu[23:16], 8'b0} * -24'h030)) + (({mcu[31:24], 8'b0} * -24'h01b)) + (({mcu[39:32], 8'b0} * 24'h01b)) + (({mcu[47:40], 8'b0} * 24'h030)) + (({mcu[55:48], 8'b0} * 24'h009)) + (({mcu[63:56], 8'b0} * -24'h029)) + (({mcu[71:64], 8'b0} * -24'h076)) + (({mcu[79:72], 8'b0} * 24'h01b)) + (({mcu[87:80], 8'b0} * 24'h08b)) + (({mcu[95:88], 8'b0} * 24'h04f)) + (({mcu[103:96], 8'b0} * -24'h04f)) + (({mcu[111:104], 8'b0} * -24'h08b)) + (({mcu[119:112], 8'b0} * -24'h01b)) + (({mcu[127:120], 8'b0} * 24'h076)) + (({mcu[135:128], 8'b0} * 24'h0b0)) + (({mcu[143:136], 8'b0} * -24'h029)) + (({mcu[151:144], 8'b0} * -24'h0d0)) + (({mcu[159:152], 8'b0} * -24'h076)) + (({mcu[167:160], 8'b0} * 24'h076)) + (({mcu[175:168], 8'b0} * 24'h0d0)) + (({mcu[183:176], 8'b0} * 24'h029)) + (({mcu[191:184], 8'b0} * -24'h0b0)) + (({mcu[199:192], 8'b0} * -24'h0d0)) + (({mcu[207:200], 8'b0} * 24'h030)) + (({mcu[215:208], 8'b0} * 24'h0f6)) + (({mcu[223:216], 8'b0} * 24'h08b)) + (({mcu[231:224], 8'b0} * -24'h08b)) + (({mcu[239:232], 8'b0} * -24'h0f6)) + (({mcu[247:240], 8'b0} * -24'h030)) + (({mcu[255:248], 8'b0} * 24'h0d0)) + (({mcu[263:256], 8'b0} * 24'h0d0)) + (({mcu[271:264], 8'b0} * -24'h030)) + (({mcu[279:272], 8'b0} * -24'h0f6)) + (({mcu[287:280], 8'b0} * -24'h08b)) + (({mcu[295:288], 8'b0} * 24'h08b)) + (({mcu[303:296], 8'b0} * 24'h0f6)) + (({mcu[311:304], 8'b0} * 24'h030)) + (({mcu[319:312], 8'b0} * -24'h0d0)) + (({mcu[327:320], 8'b0} * -24'h0b0)) + (({mcu[335:328], 8'b0} * 24'h029)) + (({mcu[343:336], 8'b0} * 24'h0d0)) + (({mcu[351:344], 8'b0} * 24'h076)) + (({mcu[359:352], 8'b0} * -24'h076)) + (({mcu[367:360], 8'b0} * -24'h0d0)) + (({mcu[375:368], 8'b0} * -24'h029)) + (({mcu[383:376], 8'b0} * 24'h0b0)) + (({mcu[391:384], 8'b0} * 24'h076)) + (({mcu[399:392], 8'b0} * -24'h01b)) + (({mcu[407:400], 8'b0} * -24'h08b)) + (({mcu[415:408], 8'b0} * -24'h04f)) + (({mcu[423:416], 8'b0} * 24'h04f)) + (({mcu[431:424], 8'b0} * 24'h08b)) + (({mcu[439:432], 8'b0} * 24'h01b)) + (({mcu[447:440], 8'b0} * -24'h076)) + (({mcu[455:448], 8'b0} * -24'h029)) + (({mcu[463:456], 8'b0} * 24'h009)) + (({mcu[471:464], 8'b0} * 24'h030)) + (({mcu[479:472], 8'b0} * 24'h01b)) + (({mcu[487:480], 8'b0} * -24'h01b)) + (({mcu[495:488], 8'b0} * -24'h030)) + (({mcu[503:496], 8'b0} * -24'h009)) + (({mcu[511:504], 8'b0} * 24'h029));
	wire[47:0] cos74_term = (({mcu[7:0], 8'b0} * 24'h023)) + (({mcu[15:8], 8'b0} * -24'h023)) + (({mcu[23:16], 8'b0} * -24'h023)) + (({mcu[31:24], 8'b0} * 24'h023)) + (({mcu[39:32], 8'b0} * 24'h023)) + (({mcu[47:40], 8'b0} * -24'h023)) + (({mcu[55:48], 8'b0} * -24'h023)) + (({mcu[63:56], 8'b0} * 24'h023)) + (({mcu[71:64], 8'b0} * -24'h064)) + (({mcu[79:72], 8'b0} * 24'h064)) + (({mcu[87:80], 8'b0} * 24'h064)) + (({mcu[95:88], 8'b0} * -24'h064)) + (({mcu[103:96], 8'b0} * -24'h064)) + (({mcu[111:104], 8'b0} * 24'h064)) + (({mcu[119:112], 8'b0} * 24'h064)) + (({mcu[127:120], 8'b0} * -24'h064)) + (({mcu[135:128], 8'b0} * 24'h096)) + (({mcu[143:136], 8'b0} * -24'h096)) + (({mcu[151:144], 8'b0} * -24'h096)) + (({mcu[159:152], 8'b0} * 24'h096)) + (({mcu[167:160], 8'b0} * 24'h096)) + (({mcu[175:168], 8'b0} * -24'h096)) + (({mcu[183:176], 8'b0} * -24'h096)) + (({mcu[191:184], 8'b0} * 24'h096)) + (({mcu[199:192], 8'b0} * -24'h0b1)) + (({mcu[207:200], 8'b0} * 24'h0b1)) + (({mcu[215:208], 8'b0} * 24'h0b1)) + (({mcu[223:216], 8'b0} * -24'h0b1)) + (({mcu[231:224], 8'b0} * -24'h0b1)) + (({mcu[239:232], 8'b0} * 24'h0b1)) + (({mcu[247:240], 8'b0} * 24'h0b1)) + (({mcu[255:248], 8'b0} * -24'h0b1)) + (({mcu[263:256], 8'b0} * 24'h0b1)) + (({mcu[271:264], 8'b0} * -24'h0b1)) + (({mcu[279:272], 8'b0} * -24'h0b1)) + (({mcu[287:280], 8'b0} * 24'h0b1)) + (({mcu[295:288], 8'b0} * 24'h0b1)) + (({mcu[303:296], 8'b0} * -24'h0b1)) + (({mcu[311:304], 8'b0} * -24'h0b1)) + (({mcu[319:312], 8'b0} * 24'h0b1)) + (({mcu[327:320], 8'b0} * -24'h096)) + (({mcu[335:328], 8'b0} * 24'h096)) + (({mcu[343:336], 8'b0} * 24'h096)) + (({mcu[351:344], 8'b0} * -24'h096)) + (({mcu[359:352], 8'b0} * -24'h096)) + (({mcu[367:360], 8'b0} * 24'h096)) + (({mcu[375:368], 8'b0} * 24'h096)) + (({mcu[383:376], 8'b0} * -24'h096)) + (({mcu[391:384], 8'b0} * 24'h064)) + (({mcu[399:392], 8'b0} * -24'h064)) + (({mcu[407:400], 8'b0} * -24'h064)) + (({mcu[415:408], 8'b0} * 24'h064)) + (({mcu[423:416], 8'b0} * 24'h064)) + (({mcu[431:424], 8'b0} * -24'h064)) + (({mcu[439:432], 8'b0} * -24'h064)) + (({mcu[447:440], 8'b0} * 24'h064)) + (({mcu[455:448], 8'b0} * -24'h023)) + (({mcu[463:456], 8'b0} * 24'h023)) + (({mcu[471:464], 8'b0} * 24'h023)) + (({mcu[479:472], 8'b0} * -24'h023)) + (({mcu[487:480], 8'b0} * -24'h023)) + (({mcu[495:488], 8'b0} * 24'h023)) + (({mcu[503:496], 8'b0} * 24'h023)) + (({mcu[511:504], 8'b0} * -24'h023));
	wire[47:0] cos75_term = (({mcu[7:0], 8'b0} * 24'h01b)) + (({mcu[15:8], 8'b0} * -24'h030)) + (({mcu[23:16], 8'b0} * 24'h009)) + (({mcu[31:24], 8'b0} * 24'h029)) + (({mcu[39:32], 8'b0} * -24'h029)) + (({mcu[47:40], 8'b0} * -24'h009)) + (({mcu[55:48], 8'b0} * 24'h030)) + (({mcu[63:56], 8'b0} * -24'h01b)) + (({mcu[71:64], 8'b0} * -24'h04f)) + (({mcu[79:72], 8'b0} * 24'h08b)) + (({mcu[87:80], 8'b0} * -24'h01b)) + (({mcu[95:88], 8'b0} * -24'h076)) + (({mcu[103:96], 8'b0} * 24'h076)) + (({mcu[111:104], 8'b0} * 24'h01b)) + (({mcu[119:112], 8'b0} * -24'h08b)) + (({mcu[127:120], 8'b0} * 24'h04f)) + (({mcu[135:128], 8'b0} * 24'h076)) + (({mcu[143:136], 8'b0} * -24'h0d0)) + (({mcu[151:144], 8'b0} * 24'h029)) + (({mcu[159:152], 8'b0} * 24'h0b0)) + (({mcu[167:160], 8'b0} * -24'h0b0)) + (({mcu[175:168], 8'b0} * -24'h029)) + (({mcu[183:176], 8'b0} * 24'h0d0)) + (({mcu[191:184], 8'b0} * -24'h076)) + (({mcu[199:192], 8'b0} * -24'h08b)) + (({mcu[207:200], 8'b0} * 24'h0f6)) + (({mcu[215:208], 8'b0} * -24'h030)) + (({mcu[223:216], 8'b0} * -24'h0d0)) + (({mcu[231:224], 8'b0} * 24'h0d0)) + (({mcu[239:232], 8'b0} * 24'h030)) + (({mcu[247:240], 8'b0} * -24'h0f6)) + (({mcu[255:248], 8'b0} * 24'h08b)) + (({mcu[263:256], 8'b0} * 24'h08b)) + (({mcu[271:264], 8'b0} * -24'h0f6)) + (({mcu[279:272], 8'b0} * 24'h030)) + (({mcu[287:280], 8'b0} * 24'h0d0)) + (({mcu[295:288], 8'b0} * -24'h0d0)) + (({mcu[303:296], 8'b0} * -24'h030)) + (({mcu[311:304], 8'b0} * 24'h0f6)) + (({mcu[319:312], 8'b0} * -24'h08b)) + (({mcu[327:320], 8'b0} * -24'h076)) + (({mcu[335:328], 8'b0} * 24'h0d0)) + (({mcu[343:336], 8'b0} * -24'h029)) + (({mcu[351:344], 8'b0} * -24'h0b0)) + (({mcu[359:352], 8'b0} * 24'h0b0)) + (({mcu[367:360], 8'b0} * 24'h029)) + (({mcu[375:368], 8'b0} * -24'h0d0)) + (({mcu[383:376], 8'b0} * 24'h076)) + (({mcu[391:384], 8'b0} * 24'h04f)) + (({mcu[399:392], 8'b0} * -24'h08b)) + (({mcu[407:400], 8'b0} * 24'h01b)) + (({mcu[415:408], 8'b0} * 24'h076)) + (({mcu[423:416], 8'b0} * -24'h076)) + (({mcu[431:424], 8'b0} * -24'h01b)) + (({mcu[439:432], 8'b0} * 24'h08b)) + (({mcu[447:440], 8'b0} * -24'h04f)) + (({mcu[455:448], 8'b0} * -24'h01b)) + (({mcu[463:456], 8'b0} * 24'h030)) + (({mcu[471:464], 8'b0} * -24'h009)) + (({mcu[479:472], 8'b0} * -24'h029)) + (({mcu[487:480], 8'b0} * 24'h029)) + (({mcu[495:488], 8'b0} * 24'h009)) + (({mcu[503:496], 8'b0} * -24'h030)) + (({mcu[511:504], 8'b0} * 24'h01b));
	wire[47:0] cos76_term = (({mcu[7:0], 8'b0} * 24'h013)) + (({mcu[15:8], 8'b0} * -24'h02e)) + (({mcu[23:16], 8'b0} * 24'h02e)) + (({mcu[31:24], 8'b0} * -24'h013)) + (({mcu[39:32], 8'b0} * -24'h013)) + (({mcu[47:40], 8'b0} * 24'h02e)) + (({mcu[55:48], 8'b0} * -24'h02e)) + (({mcu[63:56], 8'b0} * 24'h013)) + (({mcu[71:64], 8'b0} * -24'h036)) + (({mcu[79:72], 8'b0} * 24'h083)) + (({mcu[87:80], 8'b0} * -24'h083)) + (({mcu[95:88], 8'b0} * 24'h036)) + (({mcu[103:96], 8'b0} * 24'h036)) + (({mcu[111:104], 8'b0} * -24'h083)) + (({mcu[119:112], 8'b0} * 24'h083)) + (({mcu[127:120], 8'b0} * -24'h036)) + (({mcu[135:128], 8'b0} * 24'h051)) + (({mcu[143:136], 8'b0} * -24'h0c4)) + (({mcu[151:144], 8'b0} * 24'h0c4)) + (({mcu[159:152], 8'b0} * -24'h051)) + (({mcu[167:160], 8'b0} * -24'h051)) + (({mcu[175:168], 8'b0} * 24'h0c4)) + (({mcu[183:176], 8'b0} * -24'h0c4)) + (({mcu[191:184], 8'b0} * 24'h051)) + (({mcu[199:192], 8'b0} * -24'h060)) + (({mcu[207:200], 8'b0} * 24'h0e7)) + (({mcu[215:208], 8'b0} * -24'h0e7)) + (({mcu[223:216], 8'b0} * 24'h060)) + (({mcu[231:224], 8'b0} * 24'h060)) + (({mcu[239:232], 8'b0} * -24'h0e7)) + (({mcu[247:240], 8'b0} * 24'h0e7)) + (({mcu[255:248], 8'b0} * -24'h060)) + (({mcu[263:256], 8'b0} * 24'h060)) + (({mcu[271:264], 8'b0} * -24'h0e7)) + (({mcu[279:272], 8'b0} * 24'h0e7)) + (({mcu[287:280], 8'b0} * -24'h060)) + (({mcu[295:288], 8'b0} * -24'h060)) + (({mcu[303:296], 8'b0} * 24'h0e7)) + (({mcu[311:304], 8'b0} * -24'h0e7)) + (({mcu[319:312], 8'b0} * 24'h060)) + (({mcu[327:320], 8'b0} * -24'h051)) + (({mcu[335:328], 8'b0} * 24'h0c4)) + (({mcu[343:336], 8'b0} * -24'h0c4)) + (({mcu[351:344], 8'b0} * 24'h051)) + (({mcu[359:352], 8'b0} * 24'h051)) + (({mcu[367:360], 8'b0} * -24'h0c4)) + (({mcu[375:368], 8'b0} * 24'h0c4)) + (({mcu[383:376], 8'b0} * -24'h051)) + (({mcu[391:384], 8'b0} * 24'h036)) + (({mcu[399:392], 8'b0} * -24'h083)) + (({mcu[407:400], 8'b0} * 24'h083)) + (({mcu[415:408], 8'b0} * -24'h036)) + (({mcu[423:416], 8'b0} * -24'h036)) + (({mcu[431:424], 8'b0} * 24'h083)) + (({mcu[439:432], 8'b0} * -24'h083)) + (({mcu[447:440], 8'b0} * 24'h036)) + (({mcu[455:448], 8'b0} * -24'h013)) + (({mcu[463:456], 8'b0} * 24'h02e)) + (({mcu[471:464], 8'b0} * -24'h02e)) + (({mcu[479:472], 8'b0} * 24'h013)) + (({mcu[487:480], 8'b0} * 24'h013)) + (({mcu[495:488], 8'b0} * -24'h02e)) + (({mcu[503:496], 8'b0} * 24'h02e)) + (({mcu[511:504], 8'b0} * -24'h013));
	wire[47:0] cos77_term = (({mcu[7:0], 8'b0} * 24'h009)) + (({mcu[15:8], 8'b0} * -24'h01b)) + (({mcu[23:16], 8'b0} * 24'h029)) + (({mcu[31:24], 8'b0} * -24'h030)) + (({mcu[39:32], 8'b0} * 24'h030)) + (({mcu[47:40], 8'b0} * -24'h029)) + (({mcu[55:48], 8'b0} * 24'h01b)) + (({mcu[63:56], 8'b0} * -24'h009)) + (({mcu[71:64], 8'b0} * -24'h01b)) + (({mcu[79:72], 8'b0} * 24'h04f)) + (({mcu[87:80], 8'b0} * -24'h076)) + (({mcu[95:88], 8'b0} * 24'h08b)) + (({mcu[103:96], 8'b0} * -24'h08b)) + (({mcu[111:104], 8'b0} * 24'h076)) + (({mcu[119:112], 8'b0} * -24'h04f)) + (({mcu[127:120], 8'b0} * 24'h01b)) + (({mcu[135:128], 8'b0} * 24'h029)) + (({mcu[143:136], 8'b0} * -24'h076)) + (({mcu[151:144], 8'b0} * 24'h0b0)) + (({mcu[159:152], 8'b0} * -24'h0d0)) + (({mcu[167:160], 8'b0} * 24'h0d0)) + (({mcu[175:168], 8'b0} * -24'h0b0)) + (({mcu[183:176], 8'b0} * 24'h076)) + (({mcu[191:184], 8'b0} * -24'h029)) + (({mcu[199:192], 8'b0} * -24'h030)) + (({mcu[207:200], 8'b0} * 24'h08b)) + (({mcu[215:208], 8'b0} * -24'h0d0)) + (({mcu[223:216], 8'b0} * 24'h0f6)) + (({mcu[231:224], 8'b0} * -24'h0f6)) + (({mcu[239:232], 8'b0} * 24'h0d0)) + (({mcu[247:240], 8'b0} * -24'h08b)) + (({mcu[255:248], 8'b0} * 24'h030)) + (({mcu[263:256], 8'b0} * 24'h030)) + (({mcu[271:264], 8'b0} * -24'h08b)) + (({mcu[279:272], 8'b0} * 24'h0d0)) + (({mcu[287:280], 8'b0} * -24'h0f6)) + (({mcu[295:288], 8'b0} * 24'h0f6)) + (({mcu[303:296], 8'b0} * -24'h0d0)) + (({mcu[311:304], 8'b0} * 24'h08b)) + (({mcu[319:312], 8'b0} * -24'h030)) + (({mcu[327:320], 8'b0} * -24'h029)) + (({mcu[335:328], 8'b0} * 24'h076)) + (({mcu[343:336], 8'b0} * -24'h0b0)) + (({mcu[351:344], 8'b0} * 24'h0d0)) + (({mcu[359:352], 8'b0} * -24'h0d0)) + (({mcu[367:360], 8'b0} * 24'h0b0)) + (({mcu[375:368], 8'b0} * -24'h076)) + (({mcu[383:376], 8'b0} * 24'h029)) + (({mcu[391:384], 8'b0} * 24'h01b)) + (({mcu[399:392], 8'b0} * -24'h04f)) + (({mcu[407:400], 8'b0} * 24'h076)) + (({mcu[415:408], 8'b0} * -24'h08b)) + (({mcu[423:416], 8'b0} * 24'h08b)) + (({mcu[431:424], 8'b0} * -24'h076)) + (({mcu[439:432], 8'b0} * 24'h04f)) + (({mcu[447:440], 8'b0} * -24'h01b)) + (({mcu[455:448], 8'b0} * -24'h009)) + (({mcu[463:456], 8'b0} * 24'h01b)) + (({mcu[471:464], 8'b0} * -24'h029)) + (({mcu[479:472], 8'b0} * 24'h030)) + (({mcu[487:480], 8'b0} * -24'h030)) + (({mcu[495:488], 8'b0} * 24'h029)) + (({mcu[503:496], 8'b0} * -24'h01b)) + (({mcu[511:504], 8'b0} * 24'h009));

	always_comb begin
		dct[15:0] = {cos00_term, 8'b0} / 24'h10_00;
		dct[31:16] = cos01_term / 24'h0B_00;
		dct[47:32] = cos02_term[31:8] / 24'h0A_00;
		dct[63:48] = cos03_term[31:8] / 24'h10_00;
		dct[79:64] = cos04_term[31:8] / 24'h18_00;
		dct[95:80] = cos05_term[31:8] / 24'h28_00;
		dct[111:96] = cos06_term[31:8] / 24'h33_00;
		dct[127:112] = cos07_term[31:8] / 24'h3d_00;
		dct[143:128] = cos10_term[31:8] / 24'h0c_00;
		dct[159:144] = cos11_term[31:8] / 24'h0c_00;
		dct[175:160] = cos12_term[31:8] / 24'h0e_00;
		dct[191:176] = cos13_term[31:8] / 24'h13_00;
		dct[207:192] = cos14_term[31:8] / 24'h1a_00;
		dct[223:208] = cos15_term[31:8] / 24'h3a_00;
		dct[239:224] = cos16_term[31:8] / 24'h3c_00;
		dct[255:240] = cos17_term[31:8] / 24'h37_00;
		dct[271:256] = cos20_term[31:8] / 24'h0e_00;
		dct[287:272] = cos21_term[31:8] / 24'h0d_00;
		dct[303:288] = cos22_term[31:8] / 24'h10_00;
		dct[319:304] = cos23_term[31:8] / 24'h18_00;
		dct[335:320] = cos24_term[31:8] / 24'h28_00;
		dct[351:336] = cos25_term[31:8] / 24'h39_00;
		dct[367:352] = cos26_term[31:8] / 24'h45_00;
		dct[383:368] = cos27_term[31:8] / 24'h38_00;
		dct[399:384] = cos30_term[31:8] / 24'h0e_00;
		dct[415:400] = cos31_term[31:8] / 24'h11_00;
		dct[431:416] = cos32_term[31:8] / 24'h16_00;
		dct[447:432] = cos33_term[31:8] / 24'h1d_00;
		dct[463:448] = cos34_term[31:8] / 24'h33_00;
		dct[479:464] = cos35_term[31:8] / 24'h57_00;
		dct[495:480] = cos36_term[31:8] / 24'h57_00;
		dct[511:496] = cos37_term[31:8] / 24'h3e_00;
		dct[527:512] = cos40_term[31:8] / 24'h12_00;
		dct[543:528] = cos41_term[31:8] / 24'h16_00;
		dct[559:544] = cos42_term[31:8] / 24'h25_00;
		dct[575:560] = cos43_term[31:8] / 24'h38_00;
		dct[591:576] = cos44_term[31:8] / 24'h44_00;
		dct[607:592] = cos45_term[31:8] / 24'h6d_00;
		dct[623:608] = cos46_term[31:8] / 24'h67_00;
		dct[639:624] = cos47_term[31:8] / 24'h4d_00;
		dct[655:640] = cos50_term[31:8] / 24'h18_00;
		dct[671:656] = cos51_term[31:8] / 24'h23_00;
		dct[687:672] = cos52_term[31:8] / 24'h37_00;
		dct[703:688] = cos53_term[31:8] / 24'h40_00;
		dct[719:704] = cos54_term[31:8] / 24'h51_00;
		dct[735:720] = cos55_term[31:8] / 24'h68_00;
		dct[751:736] = cos56_term[31:8] / 24'h71_00;
		dct[767:752] = cos57_term[31:8] / 24'h5c_00;
		dct[783:768] = cos60_term[31:8] / 24'h31_00;
		dct[799:784] = cos61_term[31:8] / 24'h40_00;
		dct[815:800] = cos62_term[31:8] / 24'h4e_00;
		dct[831:816] = cos63_term[31:8] / 24'h57_00;
		dct[847:832] = cos64_term[31:8] / 24'h67_00;
		dct[863:848] = cos65_term[31:8] / 24'h79_00;
		dct[879:864] = cos66_term[31:8] / 24'h78_00;
		dct[895:880] = cos67_term[31:8] / 24'h65_00;
		dct[911:896] = cos70_term[31:8] / 24'h48_00;
		dct[927:912] = cos71_term[31:8] / 24'h5c_00;
		dct[943:928] = cos72_term[31:8] / 24'h5f_00;
		dct[959:944] = cos73_term[31:8] / 24'h62_00;
		dct[975:960] = cos74_term[31:8] / 24'h70_00;
		dct[991:976] = cos75_term[31:8] / 24'h64_00;
		dct[1007:992] = cos76_term[31:8] / 24'h67_00;
		dct[1023:1008] = cos77_term[31:8] / 24'h63_00;
	end
endmodule