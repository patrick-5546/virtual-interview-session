module mcu_mux_tb;
    logic [7:0][7:0][31:0] mcu_out;
    logic [7:0][7:0][31:0] mcu0;
    logic [7:0][7:0][31:0] mcu1;
    logic [10:0] x;
    
    initial begin
        mcu0[0][0] = 32'hff00;
        mcu0[0][1] = 32'h0000;
        mcu0[0][2] = 32'hff00;
        mcu0[0][3] = 32'h0000;
        mcu0[0][4] = 32'hff00;
        mcu0[0][5] = 32'h0000;
        mcu0[0][6] = 32'hff00;
        mcu0[0][7] = 32'h0000;
        mcu0[1][0] = 32'hff00;
        mcu0[1][1] = 32'h0000;
        mcu0[1][2] = 32'hff00;
        mcu0[1][3] = 32'h0000;
        mcu0[1][4] = 32'hff00;
        mcu0[1][5] = 32'h0000;
        mcu0[1][6] = 32'hff00;
        mcu0[1][7] = 32'h0000;
        mcu0[2][0] = 32'hff00;
        mcu0[2][1] = 32'h0000;
        mcu0[2][2] = 32'hff00;
        mcu0[2][3] = 32'h0000;
        mcu0[2][4] = 32'hff00;
        mcu0[2][5] = 32'h0000;
        mcu0[2][6] = 32'hff00;
        mcu0[2][7] = 32'h0000;
        mcu0[3][0] = 32'hff00;
        mcu0[3][1] = 32'h0000;
        mcu0[3][2] = 32'hff00;
        mcu0[3][3] = 32'h0000;
        mcu0[3][4] = 32'hff00;
        mcu0[3][5] = 32'h0000;
        mcu0[3][6] = 32'hff00;
        mcu0[3][7] = 32'h0000;
        mcu0[4][0] = 32'hff00;
        mcu0[4][1] = 32'h0000;
        mcu0[4][2] = 32'hff00;
        mcu0[4][3] = 32'h0000;
        mcu0[4][4] = 32'hff00;
        mcu0[4][5] = 32'h0000;
        mcu0[4][6] = 32'hff00;
        mcu0[4][7] = 32'h0000;
        mcu0[5][0] = 32'hff00;
        mcu0[5][1] = 32'h0000;
        mcu0[5][2] = 32'hff00;
        mcu0[5][3] = 32'h0000;
        mcu0[5][4] = 32'hff00;
        mcu0[5][5] = 32'h0000;
        mcu0[5][6] = 32'hff00;
        mcu0[5][7] = 32'h0000;
        mcu0[6][0] = 32'hff00;
        mcu0[6][1] = 32'h0000;
        mcu0[6][2] = 32'hff00;
        mcu0[6][3] = 32'h0000;
        mcu0[6][4] = 32'hff00;
        mcu0[6][5] = 32'h0000;
        mcu0[6][6] = 32'hff00;
        mcu0[6][7] = 32'h0000;
        mcu0[7][0] = 32'hff00;
        mcu0[7][1] = 32'h0000;
        mcu0[7][2] = 32'hff00;
        mcu0[7][3] = 32'h0000;
        mcu0[7][4] = 32'hff00;
        mcu0[7][5] = 32'h0000;
        mcu0[7][6] = 32'hff00;
        mcu0[7][7] = 32'h0000;

        mcu1[0][0] = 32'hff00;
        mcu1[0][1] = 32'hff00;
        mcu1[0][2] = 32'hff00;
        mcu1[0][3] = 32'hff00;
        mcu1[0][4] = 32'hff00;
        mcu1[0][5] = 32'hff00;
        mcu1[0][6] = 32'hff00;
        mcu1[0][7] = 32'hff00;
        mcu1[1][0] = 32'hff00;
        mcu1[1][1] = 32'hff00;
        mcu1[1][2] = 32'hff00;
        mcu1[1][3] = 32'hff00;
        mcu1[1][4] = 32'hff00;
        mcu1[1][5] = 32'hff00;
        mcu1[1][6] = 32'hff00;
        mcu1[1][7] = 32'hff00;
        mcu1[2][0] = 32'hff00;
        mcu1[2][1] = 32'hff00;
        mcu1[2][2] = 32'hff00;
        mcu1[2][3] = 32'hff00;
        mcu1[2][4] = 32'hff00;
        mcu1[2][5] = 32'hff00;
        mcu1[2][6] = 32'hff00;
        mcu1[2][7] = 32'hff00;
        mcu1[3][0] = 32'hff00;
        mcu1[3][1] = 32'hff00;
        mcu1[3][2] = 32'hff00;
        mcu1[3][3] = 32'hff00;
        mcu1[3][4] = 32'hff00;
        mcu1[3][5] = 32'hff00;
        mcu1[3][6] = 32'hff00;
        mcu1[3][7] = 32'hff00;
        mcu1[4][0] = 32'hff00;
        mcu1[4][1] = 32'hff00;
        mcu1[4][2] = 32'hff00;
        mcu1[4][3] = 32'hff00;
        mcu1[4][4] = 32'hff00;
        mcu1[4][5] = 32'hff00;
        mcu1[4][6] = 32'hff00;
        mcu1[4][7] = 32'hff00;
        mcu1[5][0] = 32'hff00;
        mcu1[5][1] = 32'hff00;
        mcu1[5][2] = 32'hff00;
        mcu1[5][3] = 32'hff00;
        mcu1[5][4] = 32'hff00;
        mcu1[5][5] = 32'hff00;
        mcu1[5][6] = 32'hff00;
        mcu1[5][7] = 32'hff00;
        mcu1[6][0] = 32'hff00;
        mcu1[6][1] = 32'hff00;
        mcu1[6][2] = 32'hff00;
        mcu1[6][3] = 32'hff00;
        mcu1[6][4] = 32'hff00;
        mcu1[6][5] = 32'hff00;
        mcu1[6][6] = 32'hff00;
        mcu1[6][7] = 32'hff00;
        mcu1[7][0] = 32'hff00;
        mcu1[7][1] = 32'hff00;
        mcu1[7][2] = 32'hff00;
        mcu1[7][3] = 32'hff00;
        mcu1[7][4] = 32'hff00;
        mcu1[7][5] = 32'hff00;
        mcu1[7][6] = 32'hff00;
        mcu1[7][7] = 32'hff00;
    end

    mcu_mux dut(.x(x), .mcu0(mcu0), .mcu1(mcu1), .mcu_out(mcu_out));
    
    initial begin
        for(int i = 208; i <= 208 + 15; i++) begin
            x = ((i - 208) / 8);
            #5;
        end
        $stop;
    end
endmodule